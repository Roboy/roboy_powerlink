// soc_system.v

// Generated using ACDS version 14.0 200 at 2018.02.08.18:45:53

`timescale 1 ps / 1 ps
module soc_system (
		input  wire        clk_50_clk,                            //                         clk_50.clk
		input  wire        reset_reset_n,                         //                          reset.reset_n
		output wire [14:0] memory_mem_a,                          //                         memory.mem_a
		output wire [2:0]  memory_mem_ba,                         //                               .mem_ba
		output wire        memory_mem_ck,                         //                               .mem_ck
		output wire        memory_mem_ck_n,                       //                               .mem_ck_n
		output wire        memory_mem_cke,                        //                               .mem_cke
		output wire        memory_mem_cs_n,                       //                               .mem_cs_n
		output wire        memory_mem_ras_n,                      //                               .mem_ras_n
		output wire        memory_mem_cas_n,                      //                               .mem_cas_n
		output wire        memory_mem_we_n,                       //                               .mem_we_n
		output wire        memory_mem_reset_n,                    //                               .mem_reset_n
		inout  wire [31:0] memory_mem_dq,                         //                               .mem_dq
		inout  wire [3:0]  memory_mem_dqs,                        //                               .mem_dqs
		inout  wire [3:0]  memory_mem_dqs_n,                      //                               .mem_dqs_n
		output wire        memory_mem_odt,                        //                               .mem_odt
		output wire [3:0]  memory_mem_dm,                         //                               .mem_dm
		input  wire        memory_oct_rzqin,                      //                               .oct_rzqin
		output wire        hps_io_hps_io_emac1_inst_TX_CLK,       //                         hps_io.hps_io_emac1_inst_TX_CLK
		output wire        hps_io_hps_io_emac1_inst_TXD0,         //                               .hps_io_emac1_inst_TXD0
		output wire        hps_io_hps_io_emac1_inst_TXD1,         //                               .hps_io_emac1_inst_TXD1
		output wire        hps_io_hps_io_emac1_inst_TXD2,         //                               .hps_io_emac1_inst_TXD2
		output wire        hps_io_hps_io_emac1_inst_TXD3,         //                               .hps_io_emac1_inst_TXD3
		input  wire        hps_io_hps_io_emac1_inst_RXD0,         //                               .hps_io_emac1_inst_RXD0
		inout  wire        hps_io_hps_io_emac1_inst_MDIO,         //                               .hps_io_emac1_inst_MDIO
		output wire        hps_io_hps_io_emac1_inst_MDC,          //                               .hps_io_emac1_inst_MDC
		input  wire        hps_io_hps_io_emac1_inst_RX_CTL,       //                               .hps_io_emac1_inst_RX_CTL
		output wire        hps_io_hps_io_emac1_inst_TX_CTL,       //                               .hps_io_emac1_inst_TX_CTL
		input  wire        hps_io_hps_io_emac1_inst_RX_CLK,       //                               .hps_io_emac1_inst_RX_CLK
		input  wire        hps_io_hps_io_emac1_inst_RXD1,         //                               .hps_io_emac1_inst_RXD1
		input  wire        hps_io_hps_io_emac1_inst_RXD2,         //                               .hps_io_emac1_inst_RXD2
		input  wire        hps_io_hps_io_emac1_inst_RXD3,         //                               .hps_io_emac1_inst_RXD3
		inout  wire        hps_io_hps_io_sdio_inst_CMD,           //                               .hps_io_sdio_inst_CMD
		inout  wire        hps_io_hps_io_sdio_inst_D0,            //                               .hps_io_sdio_inst_D0
		inout  wire        hps_io_hps_io_sdio_inst_D1,            //                               .hps_io_sdio_inst_D1
		output wire        hps_io_hps_io_sdio_inst_CLK,           //                               .hps_io_sdio_inst_CLK
		inout  wire        hps_io_hps_io_sdio_inst_D2,            //                               .hps_io_sdio_inst_D2
		inout  wire        hps_io_hps_io_sdio_inst_D3,            //                               .hps_io_sdio_inst_D3
		inout  wire        hps_io_hps_io_usb1_inst_D0,            //                               .hps_io_usb1_inst_D0
		inout  wire        hps_io_hps_io_usb1_inst_D1,            //                               .hps_io_usb1_inst_D1
		inout  wire        hps_io_hps_io_usb1_inst_D2,            //                               .hps_io_usb1_inst_D2
		inout  wire        hps_io_hps_io_usb1_inst_D3,            //                               .hps_io_usb1_inst_D3
		inout  wire        hps_io_hps_io_usb1_inst_D4,            //                               .hps_io_usb1_inst_D4
		inout  wire        hps_io_hps_io_usb1_inst_D5,            //                               .hps_io_usb1_inst_D5
		inout  wire        hps_io_hps_io_usb1_inst_D6,            //                               .hps_io_usb1_inst_D6
		inout  wire        hps_io_hps_io_usb1_inst_D7,            //                               .hps_io_usb1_inst_D7
		input  wire        hps_io_hps_io_usb1_inst_CLK,           //                               .hps_io_usb1_inst_CLK
		output wire        hps_io_hps_io_usb1_inst_STP,           //                               .hps_io_usb1_inst_STP
		input  wire        hps_io_hps_io_usb1_inst_DIR,           //                               .hps_io_usb1_inst_DIR
		input  wire        hps_io_hps_io_usb1_inst_NXT,           //                               .hps_io_usb1_inst_NXT
		output wire        hps_io_hps_io_spim1_inst_CLK,          //                               .hps_io_spim1_inst_CLK
		output wire        hps_io_hps_io_spim1_inst_MOSI,         //                               .hps_io_spim1_inst_MOSI
		input  wire        hps_io_hps_io_spim1_inst_MISO,         //                               .hps_io_spim1_inst_MISO
		output wire        hps_io_hps_io_spim1_inst_SS0,          //                               .hps_io_spim1_inst_SS0
		input  wire        hps_io_hps_io_uart0_inst_RX,           //                               .hps_io_uart0_inst_RX
		output wire        hps_io_hps_io_uart0_inst_TX,           //                               .hps_io_uart0_inst_TX
		inout  wire        hps_io_hps_io_i2c0_inst_SDA,           //                               .hps_io_i2c0_inst_SDA
		inout  wire        hps_io_hps_io_i2c0_inst_SCL,           //                               .hps_io_i2c0_inst_SCL
		inout  wire        hps_io_hps_io_i2c1_inst_SDA,           //                               .hps_io_i2c1_inst_SDA
		inout  wire        hps_io_hps_io_i2c1_inst_SCL,           //                               .hps_io_i2c1_inst_SCL
		inout  wire        hps_io_hps_io_gpio_inst_GPIO09,        //                               .hps_io_gpio_inst_GPIO09
		inout  wire        hps_io_hps_io_gpio_inst_GPIO35,        //                               .hps_io_gpio_inst_GPIO35
		inout  wire        hps_io_hps_io_gpio_inst_GPIO40,        //                               .hps_io_gpio_inst_GPIO40
		inout  wire        hps_io_hps_io_gpio_inst_GPIO53,        //                               .hps_io_gpio_inst_GPIO53
		inout  wire        hps_io_hps_io_gpio_inst_GPIO54,        //                               .hps_io_gpio_inst_GPIO54
		inout  wire        hps_io_hps_io_gpio_inst_GPIO61,        //                               .hps_io_gpio_inst_GPIO61
		input  wire        reset_1_reset_n,                       //                        reset_1.reset_n
		input  wire [3:0]  dipsw_pio_external_connection_export,  //  dipsw_pio_external_connection.export
		input  wire [1:0]  button_pio_external_connection_export, // button_pio_external_connection.export
		input  wire        hps_0_f2h_cold_reset_req_reset_n,      //       hps_0_f2h_cold_reset_req.reset_n
		input  wire        hps_0_f2h_debug_reset_req_reset_n,     //      hps_0_f2h_debug_reset_req.reset_n
		input  wire        hps_0_f2h_warm_reset_req_reset_n,      //       hps_0_f2h_warm_reset_req.reset_n
		input  wire [31:0] host_0_hps_0_h2f_gp_gp_in,             //            host_0_hps_0_h2f_gp.gp_in
		output wire [31:0] host_0_hps_0_h2f_gp_gp_out,            //                               .gp_out
		output wire        host_0_hps_0_h2f_cold_reset_reset_n,   //    host_0_hps_0_h2f_cold_reset.reset_n
		output wire [7:0]  pcp_0_benchmark_pio_export,            //            pcp_0_benchmark_pio.export
		input  wire        pcp_0_cpu_resetrequest_resetrequest,   //         pcp_0_cpu_resetrequest.resetrequest
		output wire        pcp_0_cpu_resetrequest_resettaken,     //                               .resettaken
		output wire [1:0]  powerlink_led_export,                  //                  powerlink_led.export
		output wire        openmac_0_pktactivity_export,          //          openmac_0_pktactivity.export
		output wire [0:0]  openmac_0_rmii_txEnable,               //                 openmac_0_rmii.txEnable
		output wire [1:0]  openmac_0_rmii_txData,                 //                               .txData
		input  wire [0:0]  openmac_0_rmii_rxError,                //                               .rxError
		input  wire [0:0]  openmac_0_rmii_rxCrsDataValid,         //                               .rxCrsDataValid
		input  wire [1:0]  openmac_0_rmii_rxData,                 //                               .rxData
		output wire [0:0]  openmac_0_smi_coe_smi_nPhyRst,         //                  openmac_0_smi.coe_smi_nPhyRst
		output wire [0:0]  openmac_0_smi_coe_smi_clk,             //                               .coe_smi_clk
		input  wire [0:0]  openmac_0_smi_smi_data_in,             //                               .smi_data_in
		output wire [0:0]  openmac_0_smi_smi_data_out,            //                               .smi_data_out
		output wire [0:0]  openmac_0_smi_smi_data_outEnable       //                               .smi_data_outEnable
	);

	wire         clk_100_outclk0_clk;                                 // clk_100:outclk_0 -> [host_0:clk100_clk, mm_interconnect_0:clk_100_outclk0_clk, mm_interconnect_1:clk_100_outclk0_clk, openmac_0:csi_dmaClk_clock, openmac_0:csi_mainClkx2_clock, openmac_0:csi_pktClk_clock, pcp_0:clk100_clk, rst_controller_001:clk]
	wire   [0:0] host_0_lw_bridge_m0_burstcount;                      // host_0:lw_bridge_m0_burstcount -> mm_interconnect_0:host_0_lw_bridge_m0_burstcount
	wire         host_0_lw_bridge_m0_waitrequest;                     // mm_interconnect_0:host_0_lw_bridge_m0_waitrequest -> host_0:lw_bridge_m0_waitrequest
	wire  [17:0] host_0_lw_bridge_m0_address;                         // host_0:lw_bridge_m0_address -> mm_interconnect_0:host_0_lw_bridge_m0_address
	wire  [31:0] host_0_lw_bridge_m0_writedata;                       // host_0:lw_bridge_m0_writedata -> mm_interconnect_0:host_0_lw_bridge_m0_writedata
	wire         host_0_lw_bridge_m0_write;                           // host_0:lw_bridge_m0_write -> mm_interconnect_0:host_0_lw_bridge_m0_write
	wire         host_0_lw_bridge_m0_read;                            // host_0:lw_bridge_m0_read -> mm_interconnect_0:host_0_lw_bridge_m0_read
	wire  [31:0] host_0_lw_bridge_m0_readdata;                        // mm_interconnect_0:host_0_lw_bridge_m0_readdata -> host_0:lw_bridge_m0_readdata
	wire         host_0_lw_bridge_m0_debugaccess;                     // host_0:lw_bridge_m0_debugaccess -> mm_interconnect_0:host_0_lw_bridge_m0_debugaccess
	wire   [3:0] host_0_lw_bridge_m0_byteenable;                      // host_0:lw_bridge_m0_byteenable -> mm_interconnect_0:host_0_lw_bridge_m0_byteenable
	wire         host_0_lw_bridge_m0_readdatavalid;                   // mm_interconnect_0:host_0_lw_bridge_m0_readdatavalid -> host_0:lw_bridge_m0_readdatavalid
	wire   [0:0] pcp_0_slow_bridge_burstcount;                        // pcp_0:slow_bridge_burstcount -> mm_interconnect_0:pcp_0_slow_bridge_burstcount
	wire         pcp_0_slow_bridge_waitrequest;                       // mm_interconnect_0:pcp_0_slow_bridge_waitrequest -> pcp_0:slow_bridge_waitrequest
	wire  [18:0] pcp_0_slow_bridge_address;                           // pcp_0:slow_bridge_address -> mm_interconnect_0:pcp_0_slow_bridge_address
	wire  [31:0] pcp_0_slow_bridge_writedata;                         // pcp_0:slow_bridge_writedata -> mm_interconnect_0:pcp_0_slow_bridge_writedata
	wire         pcp_0_slow_bridge_write;                             // pcp_0:slow_bridge_write -> mm_interconnect_0:pcp_0_slow_bridge_write
	wire         pcp_0_slow_bridge_read;                              // pcp_0:slow_bridge_read -> mm_interconnect_0:pcp_0_slow_bridge_read
	wire  [31:0] pcp_0_slow_bridge_readdata;                          // mm_interconnect_0:pcp_0_slow_bridge_readdata -> pcp_0:slow_bridge_readdata
	wire         pcp_0_slow_bridge_debugaccess;                       // pcp_0:slow_bridge_debugaccess -> mm_interconnect_0:pcp_0_slow_bridge_debugaccess
	wire   [3:0] pcp_0_slow_bridge_byteenable;                        // pcp_0:slow_bridge_byteenable -> mm_interconnect_0:pcp_0_slow_bridge_byteenable
	wire         pcp_0_slow_bridge_readdatavalid;                     // mm_interconnect_0:pcp_0_slow_bridge_readdatavalid -> pcp_0:slow_bridge_readdatavalid
	wire   [0:0] mm_interconnect_0_sysid_qsys_control_slave_address;  // mm_interconnect_0:sysid_qsys_control_slave_address -> sysid_qsys:address
	wire  [31:0] mm_interconnect_0_sysid_qsys_control_slave_readdata; // sysid_qsys:readdata -> mm_interconnect_0:sysid_qsys_control_slave_readdata
	wire  [31:0] mm_interconnect_0_com_mem_s1_writedata;              // mm_interconnect_0:com_mem_s1_writedata -> com_mem:writedata
	wire  [10:0] mm_interconnect_0_com_mem_s1_address;                // mm_interconnect_0:com_mem_s1_address -> com_mem:address
	wire         mm_interconnect_0_com_mem_s1_chipselect;             // mm_interconnect_0:com_mem_s1_chipselect -> com_mem:chipselect
	wire         mm_interconnect_0_com_mem_s1_clken;                  // mm_interconnect_0:com_mem_s1_clken -> com_mem:clken
	wire         mm_interconnect_0_com_mem_s1_write;                  // mm_interconnect_0:com_mem_s1_write -> com_mem:write
	wire  [31:0] mm_interconnect_0_com_mem_s1_readdata;               // com_mem:readdata -> mm_interconnect_0:com_mem_s1_readdata
	wire   [3:0] mm_interconnect_0_com_mem_s1_byteenable;             // mm_interconnect_0:com_mem_s1_byteenable -> com_mem:byteenable
	wire         mm_interconnect_0_openmac_0_macreg_waitrequest;      // openmac_0:avs_macReg_waitrequest -> mm_interconnect_0:openmac_0_macReg_waitrequest
	wire  [15:0] mm_interconnect_0_openmac_0_macreg_writedata;        // mm_interconnect_0:openmac_0_macReg_writedata -> openmac_0:avs_macReg_writedata
	wire  [11:0] mm_interconnect_0_openmac_0_macreg_address;          // mm_interconnect_0:openmac_0_macReg_address -> openmac_0:avs_macReg_address
	wire         mm_interconnect_0_openmac_0_macreg_chipselect;       // mm_interconnect_0:openmac_0_macReg_chipselect -> openmac_0:avs_macReg_chipselect
	wire         mm_interconnect_0_openmac_0_macreg_write;            // mm_interconnect_0:openmac_0_macReg_write -> openmac_0:avs_macReg_write
	wire         mm_interconnect_0_openmac_0_macreg_read;             // mm_interconnect_0:openmac_0_macReg_read -> openmac_0:avs_macReg_read
	wire  [15:0] mm_interconnect_0_openmac_0_macreg_readdata;         // openmac_0:avs_macReg_readdata -> mm_interconnect_0:openmac_0_macReg_readdata
	wire   [1:0] mm_interconnect_0_openmac_0_macreg_byteenable;       // mm_interconnect_0:openmac_0_macReg_byteenable -> openmac_0:avs_macReg_byteenable
	wire         mm_interconnect_0_openmac_0_mactimer_waitrequest;    // openmac_0:avs_macTimer_waitrequest -> mm_interconnect_0:openmac_0_macTimer_waitrequest
	wire  [31:0] mm_interconnect_0_openmac_0_mactimer_writedata;      // mm_interconnect_0:openmac_0_macTimer_writedata -> openmac_0:avs_macTimer_writedata
	wire   [2:0] mm_interconnect_0_openmac_0_mactimer_address;        // mm_interconnect_0:openmac_0_macTimer_address -> openmac_0:avs_macTimer_address
	wire         mm_interconnect_0_openmac_0_mactimer_chipselect;     // mm_interconnect_0:openmac_0_macTimer_chipselect -> openmac_0:avs_macTimer_chipselect
	wire         mm_interconnect_0_openmac_0_mactimer_write;          // mm_interconnect_0:openmac_0_macTimer_write -> openmac_0:avs_macTimer_write
	wire         mm_interconnect_0_openmac_0_mactimer_read;           // mm_interconnect_0:openmac_0_macTimer_read -> openmac_0:avs_macTimer_read
	wire  [31:0] mm_interconnect_0_openmac_0_mactimer_readdata;       // openmac_0:avs_macTimer_readdata -> mm_interconnect_0:openmac_0_macTimer_readdata
	wire   [3:0] mm_interconnect_0_openmac_0_mactimer_byteenable;     // mm_interconnect_0:openmac_0_macTimer_byteenable -> openmac_0:avs_macTimer_byteenable
	wire         mm_interconnect_0_openmac_0_pktbuf_waitrequest;      // openmac_0:avs_pktBuf_waitrequest -> mm_interconnect_0:openmac_0_pktBuf_waitrequest
	wire  [31:0] mm_interconnect_0_openmac_0_pktbuf_writedata;        // mm_interconnect_0:openmac_0_pktBuf_writedata -> openmac_0:avs_pktBuf_writedata
	wire  [12:0] mm_interconnect_0_openmac_0_pktbuf_address;          // mm_interconnect_0:openmac_0_pktBuf_address -> openmac_0:avs_pktBuf_address
	wire         mm_interconnect_0_openmac_0_pktbuf_chipselect;       // mm_interconnect_0:openmac_0_pktBuf_chipselect -> openmac_0:avs_pktBuf_chipselect
	wire         mm_interconnect_0_openmac_0_pktbuf_write;            // mm_interconnect_0:openmac_0_pktBuf_write -> openmac_0:avs_pktBuf_write
	wire         mm_interconnect_0_openmac_0_pktbuf_read;             // mm_interconnect_0:openmac_0_pktBuf_read -> openmac_0:avs_pktBuf_read
	wire  [31:0] mm_interconnect_0_openmac_0_pktbuf_readdata;         // openmac_0:avs_pktBuf_readdata -> mm_interconnect_0:openmac_0_pktBuf_readdata
	wire   [3:0] mm_interconnect_0_openmac_0_pktbuf_byteenable;       // mm_interconnect_0:openmac_0_pktBuf_byteenable -> openmac_0:avs_pktBuf_byteenable
	wire  [31:0] mm_interconnect_0_com_mem_s2_writedata;              // mm_interconnect_0:com_mem_s2_writedata -> com_mem:writedata2
	wire  [10:0] mm_interconnect_0_com_mem_s2_address;                // mm_interconnect_0:com_mem_s2_address -> com_mem:address2
	wire         mm_interconnect_0_com_mem_s2_chipselect;             // mm_interconnect_0:com_mem_s2_chipselect -> com_mem:chipselect2
	wire         mm_interconnect_0_com_mem_s2_clken;                  // mm_interconnect_0:com_mem_s2_clken -> com_mem:clken2
	wire         mm_interconnect_0_com_mem_s2_write;                  // mm_interconnect_0:com_mem_s2_write -> com_mem:write2
	wire  [31:0] mm_interconnect_0_com_mem_s2_readdata;               // com_mem:readdata2 -> mm_interconnect_0:com_mem_s2_readdata
	wire   [3:0] mm_interconnect_0_com_mem_s2_byteenable;             // mm_interconnect_0:com_mem_s2_byteenable -> com_mem:byteenable2
	wire  [12:0] openmac_0_dma_burstcount;                            // openmac_0:avm_dma_burstcount -> mm_interconnect_1:openmac_0_dma_burstcount
	wire         openmac_0_dma_waitrequest;                           // mm_interconnect_1:openmac_0_dma_waitrequest -> openmac_0:avm_dma_waitrequest
	wire  [15:0] openmac_0_dma_writedata;                             // openmac_0:avm_dma_writedata -> mm_interconnect_1:openmac_0_dma_writedata
	wire  [18:0] openmac_0_dma_address;                               // openmac_0:avm_dma_address -> mm_interconnect_1:openmac_0_dma_address
	wire         openmac_0_dma_write;                                 // openmac_0:avm_dma_write -> mm_interconnect_1:openmac_0_dma_write
	wire   [1:0] openmac_0_dma_byteenable;                            // openmac_0:avm_dma_byteenable -> mm_interconnect_1:openmac_0_dma_byteenable
	wire   [0:0] host_0_fpga_mem_burstcount;                          // host_0:fpga_mem_burstcount -> mm_interconnect_1:host_0_fpga_mem_burstcount
	wire         host_0_fpga_mem_waitrequest;                         // mm_interconnect_1:host_0_fpga_mem_waitrequest -> host_0:fpga_mem_waitrequest
	wire  [26:0] host_0_fpga_mem_address;                             // host_0:fpga_mem_address -> mm_interconnect_1:host_0_fpga_mem_address
	wire  [31:0] host_0_fpga_mem_writedata;                           // host_0:fpga_mem_writedata -> mm_interconnect_1:host_0_fpga_mem_writedata
	wire         host_0_fpga_mem_write;                               // host_0:fpga_mem_write -> mm_interconnect_1:host_0_fpga_mem_write
	wire         host_0_fpga_mem_read;                                // host_0:fpga_mem_read -> mm_interconnect_1:host_0_fpga_mem_read
	wire  [31:0] host_0_fpga_mem_readdata;                            // mm_interconnect_1:host_0_fpga_mem_readdata -> host_0:fpga_mem_readdata
	wire         host_0_fpga_mem_debugaccess;                         // host_0:fpga_mem_debugaccess -> mm_interconnect_1:host_0_fpga_mem_debugaccess
	wire   [3:0] host_0_fpga_mem_byteenable;                          // host_0:fpga_mem_byteenable -> mm_interconnect_1:host_0_fpga_mem_byteenable
	wire         host_0_fpga_mem_readdatavalid;                       // mm_interconnect_1:host_0_fpga_mem_readdatavalid -> host_0:fpga_mem_readdatavalid
	wire   [0:0] pcp_0_cpu_bridge_burstcount;                         // pcp_0:cpu_bridge_burstcount -> mm_interconnect_1:pcp_0_cpu_bridge_burstcount
	wire         pcp_0_cpu_bridge_waitrequest;                        // mm_interconnect_1:pcp_0_cpu_bridge_waitrequest -> pcp_0:cpu_bridge_waitrequest
	wire  [21:0] pcp_0_cpu_bridge_address;                            // pcp_0:cpu_bridge_address -> mm_interconnect_1:pcp_0_cpu_bridge_address
	wire  [31:0] pcp_0_cpu_bridge_writedata;                          // pcp_0:cpu_bridge_writedata -> mm_interconnect_1:pcp_0_cpu_bridge_writedata
	wire         pcp_0_cpu_bridge_write;                              // pcp_0:cpu_bridge_write -> mm_interconnect_1:pcp_0_cpu_bridge_write
	wire         pcp_0_cpu_bridge_read;                               // pcp_0:cpu_bridge_read -> mm_interconnect_1:pcp_0_cpu_bridge_read
	wire  [31:0] pcp_0_cpu_bridge_readdata;                           // mm_interconnect_1:pcp_0_cpu_bridge_readdata -> pcp_0:cpu_bridge_readdata
	wire         pcp_0_cpu_bridge_debugaccess;                        // pcp_0:cpu_bridge_debugaccess -> mm_interconnect_1:pcp_0_cpu_bridge_debugaccess
	wire   [3:0] pcp_0_cpu_bridge_byteenable;                         // pcp_0:cpu_bridge_byteenable -> mm_interconnect_1:pcp_0_cpu_bridge_byteenable
	wire         pcp_0_cpu_bridge_readdatavalid;                      // mm_interconnect_1:pcp_0_cpu_bridge_readdatavalid -> pcp_0:cpu_bridge_readdatavalid
	wire   [0:0] pcp_0_flash_bridge_burstcount;                       // pcp_0:flash_bridge_burstcount -> mm_interconnect_1:pcp_0_flash_bridge_burstcount
	wire         pcp_0_flash_bridge_waitrequest;                      // mm_interconnect_1:pcp_0_flash_bridge_waitrequest -> pcp_0:flash_bridge_waitrequest
	wire  [21:0] pcp_0_flash_bridge_address;                          // pcp_0:flash_bridge_address -> mm_interconnect_1:pcp_0_flash_bridge_address
	wire  [31:0] pcp_0_flash_bridge_writedata;                        // pcp_0:flash_bridge_writedata -> mm_interconnect_1:pcp_0_flash_bridge_writedata
	wire         pcp_0_flash_bridge_write;                            // pcp_0:flash_bridge_write -> mm_interconnect_1:pcp_0_flash_bridge_write
	wire         pcp_0_flash_bridge_read;                             // pcp_0:flash_bridge_read -> mm_interconnect_1:pcp_0_flash_bridge_read
	wire  [31:0] pcp_0_flash_bridge_readdata;                         // mm_interconnect_1:pcp_0_flash_bridge_readdata -> pcp_0:flash_bridge_readdata
	wire         pcp_0_flash_bridge_debugaccess;                      // pcp_0:flash_bridge_debugaccess -> mm_interconnect_1:pcp_0_flash_bridge_debugaccess
	wire   [3:0] pcp_0_flash_bridge_byteenable;                       // pcp_0:flash_bridge_byteenable -> mm_interconnect_1:pcp_0_flash_bridge_byteenable
	wire         pcp_0_flash_bridge_readdatavalid;                    // mm_interconnect_1:pcp_0_flash_bridge_readdatavalid -> pcp_0:flash_bridge_readdatavalid
	wire  [31:0] mm_interconnect_1_onchip_memory2_0_s1_writedata;     // mm_interconnect_1:onchip_memory2_0_s1_writedata -> onchip_memory2_0:writedata
	wire  [16:0] mm_interconnect_1_onchip_memory2_0_s1_address;       // mm_interconnect_1:onchip_memory2_0_s1_address -> onchip_memory2_0:address
	wire         mm_interconnect_1_onchip_memory2_0_s1_chipselect;    // mm_interconnect_1:onchip_memory2_0_s1_chipselect -> onchip_memory2_0:chipselect
	wire         mm_interconnect_1_onchip_memory2_0_s1_clken;         // mm_interconnect_1:onchip_memory2_0_s1_clken -> onchip_memory2_0:clken
	wire         mm_interconnect_1_onchip_memory2_0_s1_write;         // mm_interconnect_1:onchip_memory2_0_s1_write -> onchip_memory2_0:write
	wire  [31:0] mm_interconnect_1_onchip_memory2_0_s1_readdata;      // onchip_memory2_0:readdata -> mm_interconnect_1:onchip_memory2_0_s1_readdata
	wire   [3:0] mm_interconnect_1_onchip_memory2_0_s1_byteenable;    // mm_interconnect_1:onchip_memory2_0_s1_byteenable -> onchip_memory2_0:byteenable
	wire         irq_mapper_receiver0_irq;                            // openmac_0:ins_timerPulse_irq -> irq_mapper:receiver0_irq
	wire   [0:0] host_0_hostif_irq_i_irq;                             // irq_mapper:sender_irq -> host_0:hostif_irq_i_irq
	wire         irq_mapper_001_receiver0_irq;                        // openmac_0:ins_timerIrq_irq -> irq_mapper_001:receiver0_irq
	wire   [0:0] pcp_0_sync_irq_irq;                                  // irq_mapper_001:sender_irq -> pcp_0:sync_irq_irq
	wire         irq_mapper_002_receiver0_irq;                        // openmac_0:ins_macIrq_irq -> irq_mapper_002:receiver0_irq
	wire   [0:0] pcp_0_mac_irq_irq;                                   // irq_mapper_002:sender_irq -> pcp_0:mac_irq_irq
	wire   [3:0] pcp_0_gp_irq_irq;                                    // irq_mapper_003:sender_irq -> pcp_0:gp_irq_irq
	wire         rst_controller_reset_out_reset;                      // rst_controller:reset_out -> [clk_100:rst, com_mem:reset, com_mem:reset2, irq_mapper_001:reset, irq_mapper_002:reset, irq_mapper_003:reset, mm_interconnect_0:host_0_reset_clk50_reset_bridge_in_reset_reset, mm_interconnect_0:sysid_qsys_reset_reset_bridge_in_reset_reset, mm_interconnect_1:onchip_memory2_0_reset1_reset_bridge_in_reset_reset, onchip_memory2_0:reset, rst_translator:in_reset, sysid_qsys:reset_n]
	wire         rst_controller_reset_out_reset_req;                  // rst_controller:reset_req -> [com_mem:reset_req, com_mem:reset_req2, onchip_memory2_0:reset_req, rst_translator:reset_req_in]
	wire         rst_controller_001_reset_out_reset;                  // rst_controller_001:reset_out -> [mm_interconnect_0:openmac_0_pktBuf_translator_reset_reset_bridge_in_reset_reset, mm_interconnect_0:openmac_0_pktRst_reset_bridge_in_reset_reset, mm_interconnect_1:openmac_0_dmaRst_reset_bridge_in_reset_reset, mm_interconnect_1:openmac_0_dma_translator_reset_reset_bridge_in_reset_reset]

	soc_system_sysid_qsys sysid_qsys (
		.clock    (clk_50_clk),                                          //           clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                     //         reset.reset_n
		.readdata (mm_interconnect_0_sysid_qsys_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_sysid_qsys_control_slave_address)   //              .address
	);

	alteraOpenmacTop #(
		.gPhyPortCount          (1),
		.gPhyPortType           (1),
		.gSmiPortCount          (1),
		.gEndianness            ("little"),
		.gEnableActivity        (1),
		.gEnableDmaObserver     (1),
		.gDmaAddrWidth          (19),
		.gDmaDataWidth          (16),
		.gDmaBurstCountWidth    (13),
		.gDmaWriteBurstLength   (4),
		.gDmaReadBurstLength    (1),
		.gDmaWriteFifoLength    (16),
		.gDmaReadFifoLength     (16),
		.gPacketBufferLocTx     (1),
		.gPacketBufferLocRx     (2),
		.gPacketBufferLog2Size  (15),
		.gTimerEnablePulse      (1),
		.gTimerEnablePulseWidth (0),
		.gTimerPulseRegWidth    (10)
	) openmac_0 (
		.csi_mainClk_clock        (clk_50_clk),                                       //     mainClk.clk
		.csi_mainClkx2_clock      (clk_100_outclk0_clk),                              //   mainClkx2.clk
		.csi_dmaClk_clock         (clk_100_outclk0_clk),                              //      dmaClk.clk
		.csi_pktClk_clock         (clk_100_outclk0_clk),                              //      pktClk.clk
		.rsi_mainRst_reset        (~reset_reset_n),                                   //     mainRst.reset
		.rsi_dmaRst_reset         (~reset_reset_n),                                   //      dmaRst.reset
		.rsi_pktRst_reset         (~reset_reset_n),                                   //      pktRst.reset
		.avs_macReg_chipselect    (mm_interconnect_0_openmac_0_macreg_chipselect),    //      macReg.chipselect
		.avs_macReg_write         (mm_interconnect_0_openmac_0_macreg_write),         //            .write
		.avs_macReg_read          (mm_interconnect_0_openmac_0_macreg_read),          //            .read
		.avs_macReg_waitrequest   (mm_interconnect_0_openmac_0_macreg_waitrequest),   //            .waitrequest
		.avs_macReg_byteenable    (mm_interconnect_0_openmac_0_macreg_byteenable),    //            .byteenable
		.avs_macReg_address       (mm_interconnect_0_openmac_0_macreg_address),       //            .address
		.avs_macReg_writedata     (mm_interconnect_0_openmac_0_macreg_writedata),     //            .writedata
		.avs_macReg_readdata      (mm_interconnect_0_openmac_0_macreg_readdata),      //            .readdata
		.avs_macTimer_chipselect  (mm_interconnect_0_openmac_0_mactimer_chipselect),  //    macTimer.chipselect
		.avs_macTimer_write       (mm_interconnect_0_openmac_0_mactimer_write),       //            .write
		.avs_macTimer_read        (mm_interconnect_0_openmac_0_mactimer_read),        //            .read
		.avs_macTimer_waitrequest (mm_interconnect_0_openmac_0_mactimer_waitrequest), //            .waitrequest
		.avs_macTimer_address     (mm_interconnect_0_openmac_0_mactimer_address),     //            .address
		.avs_macTimer_byteenable  (mm_interconnect_0_openmac_0_mactimer_byteenable),  //            .byteenable
		.avs_macTimer_writedata   (mm_interconnect_0_openmac_0_mactimer_writedata),   //            .writedata
		.avs_macTimer_readdata    (mm_interconnect_0_openmac_0_mactimer_readdata),    //            .readdata
		.avs_pktBuf_chipselect    (mm_interconnect_0_openmac_0_pktbuf_chipselect),    //      pktBuf.chipselect
		.avs_pktBuf_write         (mm_interconnect_0_openmac_0_pktbuf_write),         //            .write
		.avs_pktBuf_read          (mm_interconnect_0_openmac_0_pktbuf_read),          //            .read
		.avs_pktBuf_waitrequest   (mm_interconnect_0_openmac_0_pktbuf_waitrequest),   //            .waitrequest
		.avs_pktBuf_byteenable    (mm_interconnect_0_openmac_0_pktbuf_byteenable),    //            .byteenable
		.avs_pktBuf_address       (mm_interconnect_0_openmac_0_pktbuf_address),       //            .address
		.avs_pktBuf_writedata     (mm_interconnect_0_openmac_0_pktbuf_writedata),     //            .writedata
		.avs_pktBuf_readdata      (mm_interconnect_0_openmac_0_pktbuf_readdata),      //            .readdata
		.avm_dma_write            (openmac_0_dma_write),                              //         dma.write
		.avm_dma_waitrequest      (openmac_0_dma_waitrequest),                        //            .waitrequest
		.avm_dma_byteenable       (openmac_0_dma_byteenable),                         //            .byteenable
		.avm_dma_address          (openmac_0_dma_address),                            //            .address
		.avm_dma_burstcount       (openmac_0_dma_burstcount),                         //            .burstcount
		.avm_dma_writedata        (openmac_0_dma_writedata),                          //            .writedata
		.ins_timerIrq_irq         (irq_mapper_001_receiver0_irq),                     //    timerIrq.irq
		.ins_timerPulse_irq       (irq_mapper_receiver0_irq),                         //  timerPulse.irq
		.ins_macIrq_irq           (irq_mapper_002_receiver0_irq),                     //      macIrq.irq
		.coe_rmii_txEnable        (openmac_0_rmii_txEnable),                          //        rmii.export
		.coe_rmii_txData          (openmac_0_rmii_txData),                            //            .export
		.coe_rmii_rxError         (openmac_0_rmii_rxError),                           //            .export
		.coe_rmii_rxCrsDataValid  (openmac_0_rmii_rxCrsDataValid),                    //            .export
		.coe_rmii_rxData          (openmac_0_rmii_rxData),                            //            .export
		.coe_smi_nPhyRst          (openmac_0_smi_coe_smi_nPhyRst),                    //         smi.export
		.coe_smi_clk              (openmac_0_smi_coe_smi_clk),                        //            .export
		.smi_data_in              (openmac_0_smi_smi_data_in),                        //            .export
		.smi_data_out             (openmac_0_smi_smi_data_out),                       //            .export
		.smi_data_outEnable       (openmac_0_smi_smi_data_outEnable),                 //            .export
		.coe_pktActivity          (openmac_0_pktactivity_export),                     // pktActivity.export
		.avm_dma_read             (),                                                 // (terminated)
		.avm_dma_readdatavalid    (1'b0),                                             // (terminated)
		.avm_dma_readdata         (16'b0000000000000000),                             // (terminated)
		.coe_mii_txEnable         (),                                                 // (terminated)
		.coe_mii_txData           (),                                                 // (terminated)
		.coe_mii_txClk            (1'b0),                                             // (terminated)
		.coe_mii_rxError          (1'b0),                                             // (terminated)
		.coe_mii_rxDataValid      (1'b0),                                             // (terminated)
		.coe_mii_rxData           (4'b0000),                                          // (terminated)
		.coe_mii_rxClk            (1'b0)                                              // (terminated)
	);

	soc_system_com_mem com_mem (
		.clk         (clk_50_clk),                              //   clk1.clk
		.address     (mm_interconnect_0_com_mem_s1_address),    //     s1.address
		.clken       (mm_interconnect_0_com_mem_s1_clken),      //       .clken
		.chipselect  (mm_interconnect_0_com_mem_s1_chipselect), //       .chipselect
		.write       (mm_interconnect_0_com_mem_s1_write),      //       .write
		.readdata    (mm_interconnect_0_com_mem_s1_readdata),   //       .readdata
		.writedata   (mm_interconnect_0_com_mem_s1_writedata),  //       .writedata
		.byteenable  (mm_interconnect_0_com_mem_s1_byteenable), //       .byteenable
		.reset       (rst_controller_reset_out_reset),          // reset1.reset
		.reset_req   (rst_controller_reset_out_reset_req),      //       .reset_req
		.address2    (mm_interconnect_0_com_mem_s2_address),    //     s2.address
		.chipselect2 (mm_interconnect_0_com_mem_s2_chipselect), //       .chipselect
		.clken2      (mm_interconnect_0_com_mem_s2_clken),      //       .clken
		.write2      (mm_interconnect_0_com_mem_s2_write),      //       .write
		.readdata2   (mm_interconnect_0_com_mem_s2_readdata),   //       .readdata
		.writedata2  (mm_interconnect_0_com_mem_s2_writedata),  //       .writedata
		.byteenable2 (mm_interconnect_0_com_mem_s2_byteenable), //       .byteenable
		.clk2        (clk_50_clk),                              //   clk2.clk
		.reset2      (rst_controller_reset_out_reset),          // reset2.reset
		.reset_req2  (rst_controller_reset_out_reset_req)       //       .reset_req
	);

	soc_system_clk_100 clk_100 (
		.refclk   (clk_50_clk),                     //  refclk.clk
		.rst      (rst_controller_reset_out_reset), //   reset.reset
		.outclk_0 (clk_100_outclk0_clk),            // outclk0.clk
		.locked   ()                                // (terminated)
	);

	soc_system_onchip_memory2_0 onchip_memory2_0 (
		.clk        (clk_50_clk),                                       //   clk1.clk
		.address    (mm_interconnect_1_onchip_memory2_0_s1_address),    //     s1.address
		.clken      (mm_interconnect_1_onchip_memory2_0_s1_clken),      //       .clken
		.chipselect (mm_interconnect_1_onchip_memory2_0_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_1_onchip_memory2_0_s1_write),      //       .write
		.readdata   (mm_interconnect_1_onchip_memory2_0_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_1_onchip_memory2_0_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_1_onchip_memory2_0_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),                   // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req)                //       .reset_req
	);

	soc_system_host_0 host_0 (
		.memory_mem_a                          (memory_mem_a),                          //                         memory.mem_a
		.memory_mem_ba                         (memory_mem_ba),                         //                               .mem_ba
		.memory_mem_ck                         (memory_mem_ck),                         //                               .mem_ck
		.memory_mem_ck_n                       (memory_mem_ck_n),                       //                               .mem_ck_n
		.memory_mem_cke                        (memory_mem_cke),                        //                               .mem_cke
		.memory_mem_cs_n                       (memory_mem_cs_n),                       //                               .mem_cs_n
		.memory_mem_ras_n                      (memory_mem_ras_n),                      //                               .mem_ras_n
		.memory_mem_cas_n                      (memory_mem_cas_n),                      //                               .mem_cas_n
		.memory_mem_we_n                       (memory_mem_we_n),                       //                               .mem_we_n
		.memory_mem_reset_n                    (memory_mem_reset_n),                    //                               .mem_reset_n
		.memory_mem_dq                         (memory_mem_dq),                         //                               .mem_dq
		.memory_mem_dqs                        (memory_mem_dqs),                        //                               .mem_dqs
		.memory_mem_dqs_n                      (memory_mem_dqs_n),                      //                               .mem_dqs_n
		.memory_mem_odt                        (memory_mem_odt),                        //                               .mem_odt
		.memory_mem_dm                         (memory_mem_dm),                         //                               .mem_dm
		.memory_oct_rzqin                      (memory_oct_rzqin),                      //                               .oct_rzqin
		.clk50_clk                             (clk_50_clk),                            //                          clk50.clk
		.reset_clk50_reset_n                   (reset_reset_n),                         //                    reset_clk50.reset_n
		.hps_0_hps_io_hps_io_emac1_inst_TX_CLK (hps_io_hps_io_emac1_inst_TX_CLK),       //                   hps_0_hps_io.hps_io_emac1_inst_TX_CLK
		.hps_0_hps_io_hps_io_emac1_inst_TXD0   (hps_io_hps_io_emac1_inst_TXD0),         //                               .hps_io_emac1_inst_TXD0
		.hps_0_hps_io_hps_io_emac1_inst_TXD1   (hps_io_hps_io_emac1_inst_TXD1),         //                               .hps_io_emac1_inst_TXD1
		.hps_0_hps_io_hps_io_emac1_inst_TXD2   (hps_io_hps_io_emac1_inst_TXD2),         //                               .hps_io_emac1_inst_TXD2
		.hps_0_hps_io_hps_io_emac1_inst_TXD3   (hps_io_hps_io_emac1_inst_TXD3),         //                               .hps_io_emac1_inst_TXD3
		.hps_0_hps_io_hps_io_emac1_inst_RXD0   (hps_io_hps_io_emac1_inst_RXD0),         //                               .hps_io_emac1_inst_RXD0
		.hps_0_hps_io_hps_io_emac1_inst_MDIO   (hps_io_hps_io_emac1_inst_MDIO),         //                               .hps_io_emac1_inst_MDIO
		.hps_0_hps_io_hps_io_emac1_inst_MDC    (hps_io_hps_io_emac1_inst_MDC),          //                               .hps_io_emac1_inst_MDC
		.hps_0_hps_io_hps_io_emac1_inst_RX_CTL (hps_io_hps_io_emac1_inst_RX_CTL),       //                               .hps_io_emac1_inst_RX_CTL
		.hps_0_hps_io_hps_io_emac1_inst_TX_CTL (hps_io_hps_io_emac1_inst_TX_CTL),       //                               .hps_io_emac1_inst_TX_CTL
		.hps_0_hps_io_hps_io_emac1_inst_RX_CLK (hps_io_hps_io_emac1_inst_RX_CLK),       //                               .hps_io_emac1_inst_RX_CLK
		.hps_0_hps_io_hps_io_emac1_inst_RXD1   (hps_io_hps_io_emac1_inst_RXD1),         //                               .hps_io_emac1_inst_RXD1
		.hps_0_hps_io_hps_io_emac1_inst_RXD2   (hps_io_hps_io_emac1_inst_RXD2),         //                               .hps_io_emac1_inst_RXD2
		.hps_0_hps_io_hps_io_emac1_inst_RXD3   (hps_io_hps_io_emac1_inst_RXD3),         //                               .hps_io_emac1_inst_RXD3
		.hps_0_hps_io_hps_io_sdio_inst_CMD     (hps_io_hps_io_sdio_inst_CMD),           //                               .hps_io_sdio_inst_CMD
		.hps_0_hps_io_hps_io_sdio_inst_D0      (hps_io_hps_io_sdio_inst_D0),            //                               .hps_io_sdio_inst_D0
		.hps_0_hps_io_hps_io_sdio_inst_D1      (hps_io_hps_io_sdio_inst_D1),            //                               .hps_io_sdio_inst_D1
		.hps_0_hps_io_hps_io_sdio_inst_CLK     (hps_io_hps_io_sdio_inst_CLK),           //                               .hps_io_sdio_inst_CLK
		.hps_0_hps_io_hps_io_sdio_inst_D2      (hps_io_hps_io_sdio_inst_D2),            //                               .hps_io_sdio_inst_D2
		.hps_0_hps_io_hps_io_sdio_inst_D3      (hps_io_hps_io_sdio_inst_D3),            //                               .hps_io_sdio_inst_D3
		.hps_0_hps_io_hps_io_usb1_inst_D0      (hps_io_hps_io_usb1_inst_D0),            //                               .hps_io_usb1_inst_D0
		.hps_0_hps_io_hps_io_usb1_inst_D1      (hps_io_hps_io_usb1_inst_D1),            //                               .hps_io_usb1_inst_D1
		.hps_0_hps_io_hps_io_usb1_inst_D2      (hps_io_hps_io_usb1_inst_D2),            //                               .hps_io_usb1_inst_D2
		.hps_0_hps_io_hps_io_usb1_inst_D3      (hps_io_hps_io_usb1_inst_D3),            //                               .hps_io_usb1_inst_D3
		.hps_0_hps_io_hps_io_usb1_inst_D4      (hps_io_hps_io_usb1_inst_D4),            //                               .hps_io_usb1_inst_D4
		.hps_0_hps_io_hps_io_usb1_inst_D5      (hps_io_hps_io_usb1_inst_D5),            //                               .hps_io_usb1_inst_D5
		.hps_0_hps_io_hps_io_usb1_inst_D6      (hps_io_hps_io_usb1_inst_D6),            //                               .hps_io_usb1_inst_D6
		.hps_0_hps_io_hps_io_usb1_inst_D7      (hps_io_hps_io_usb1_inst_D7),            //                               .hps_io_usb1_inst_D7
		.hps_0_hps_io_hps_io_usb1_inst_CLK     (hps_io_hps_io_usb1_inst_CLK),           //                               .hps_io_usb1_inst_CLK
		.hps_0_hps_io_hps_io_usb1_inst_STP     (hps_io_hps_io_usb1_inst_STP),           //                               .hps_io_usb1_inst_STP
		.hps_0_hps_io_hps_io_usb1_inst_DIR     (hps_io_hps_io_usb1_inst_DIR),           //                               .hps_io_usb1_inst_DIR
		.hps_0_hps_io_hps_io_usb1_inst_NXT     (hps_io_hps_io_usb1_inst_NXT),           //                               .hps_io_usb1_inst_NXT
		.hps_0_hps_io_hps_io_spim1_inst_CLK    (hps_io_hps_io_spim1_inst_CLK),          //                               .hps_io_spim1_inst_CLK
		.hps_0_hps_io_hps_io_spim1_inst_MOSI   (hps_io_hps_io_spim1_inst_MOSI),         //                               .hps_io_spim1_inst_MOSI
		.hps_0_hps_io_hps_io_spim1_inst_MISO   (hps_io_hps_io_spim1_inst_MISO),         //                               .hps_io_spim1_inst_MISO
		.hps_0_hps_io_hps_io_spim1_inst_SS0    (hps_io_hps_io_spim1_inst_SS0),          //                               .hps_io_spim1_inst_SS0
		.hps_0_hps_io_hps_io_uart0_inst_RX     (hps_io_hps_io_uart0_inst_RX),           //                               .hps_io_uart0_inst_RX
		.hps_0_hps_io_hps_io_uart0_inst_TX     (hps_io_hps_io_uart0_inst_TX),           //                               .hps_io_uart0_inst_TX
		.hps_0_hps_io_hps_io_i2c0_inst_SDA     (hps_io_hps_io_i2c0_inst_SDA),           //                               .hps_io_i2c0_inst_SDA
		.hps_0_hps_io_hps_io_i2c0_inst_SCL     (hps_io_hps_io_i2c0_inst_SCL),           //                               .hps_io_i2c0_inst_SCL
		.hps_0_hps_io_hps_io_i2c1_inst_SDA     (hps_io_hps_io_i2c1_inst_SDA),           //                               .hps_io_i2c1_inst_SDA
		.hps_0_hps_io_hps_io_i2c1_inst_SCL     (hps_io_hps_io_i2c1_inst_SCL),           //                               .hps_io_i2c1_inst_SCL
		.hps_0_hps_io_hps_io_gpio_inst_GPIO09  (hps_io_hps_io_gpio_inst_GPIO09),        //                               .hps_io_gpio_inst_GPIO09
		.hps_0_hps_io_hps_io_gpio_inst_GPIO35  (hps_io_hps_io_gpio_inst_GPIO35),        //                               .hps_io_gpio_inst_GPIO35
		.hps_0_hps_io_hps_io_gpio_inst_GPIO40  (hps_io_hps_io_gpio_inst_GPIO40),        //                               .hps_io_gpio_inst_GPIO40
		.hps_0_hps_io_hps_io_gpio_inst_GPIO53  (hps_io_hps_io_gpio_inst_GPIO53),        //                               .hps_io_gpio_inst_GPIO53
		.hps_0_hps_io_hps_io_gpio_inst_GPIO54  (hps_io_hps_io_gpio_inst_GPIO54),        //                               .hps_io_gpio_inst_GPIO54
		.hps_0_hps_io_hps_io_gpio_inst_GPIO61  (hps_io_hps_io_gpio_inst_GPIO61),        //                               .hps_io_gpio_inst_GPIO61
		.dipsw_pio_external_connection_export  (dipsw_pio_external_connection_export),  //  dipsw_pio_external_connection.export
		.button_pio_external_connection_export (button_pio_external_connection_export), // button_pio_external_connection.export
		.hps_0_f2h_cold_reset_req_reset_n      (hps_0_f2h_cold_reset_req_reset_n),      //       hps_0_f2h_cold_reset_req.reset_n
		.hps_0_f2h_debug_reset_req_reset_n     (hps_0_f2h_debug_reset_req_reset_n),     //      hps_0_f2h_debug_reset_req.reset_n
		.hps_0_f2h_warm_reset_req_reset_n      (hps_0_f2h_warm_reset_req_reset_n),      //       hps_0_f2h_warm_reset_req.reset_n
		.clk100_clk                            (clk_100_outclk0_clk),                   //                         clk100.clk
		.fpga_mem_waitrequest                  (host_0_fpga_mem_waitrequest),           //                       fpga_mem.waitrequest
		.fpga_mem_readdata                     (host_0_fpga_mem_readdata),              //                               .readdata
		.fpga_mem_readdatavalid                (host_0_fpga_mem_readdatavalid),         //                               .readdatavalid
		.fpga_mem_burstcount                   (host_0_fpga_mem_burstcount),            //                               .burstcount
		.fpga_mem_writedata                    (host_0_fpga_mem_writedata),             //                               .writedata
		.fpga_mem_address                      (host_0_fpga_mem_address),               //                               .address
		.fpga_mem_write                        (host_0_fpga_mem_write),                 //                               .write
		.fpga_mem_read                         (host_0_fpga_mem_read),                  //                               .read
		.fpga_mem_byteenable                   (host_0_fpga_mem_byteenable),            //                               .byteenable
		.fpga_mem_debugaccess                  (host_0_fpga_mem_debugaccess),           //                               .debugaccess
		.reset_clk100_reset_n                  (reset_1_reset_n),                       //                   reset_clk100.reset_n
		.hostif_irq_i_irq                      (host_0_hostif_irq_i_irq),               //                   hostif_irq_i.irq
		.lw_bridge_m0_waitrequest              (host_0_lw_bridge_m0_waitrequest),       //                   lw_bridge_m0.waitrequest
		.lw_bridge_m0_readdata                 (host_0_lw_bridge_m0_readdata),          //                               .readdata
		.lw_bridge_m0_readdatavalid            (host_0_lw_bridge_m0_readdatavalid),     //                               .readdatavalid
		.lw_bridge_m0_burstcount               (host_0_lw_bridge_m0_burstcount),        //                               .burstcount
		.lw_bridge_m0_writedata                (host_0_lw_bridge_m0_writedata),         //                               .writedata
		.lw_bridge_m0_address                  (host_0_lw_bridge_m0_address),           //                               .address
		.lw_bridge_m0_write                    (host_0_lw_bridge_m0_write),             //                               .write
		.lw_bridge_m0_read                     (host_0_lw_bridge_m0_read),              //                               .read
		.lw_bridge_m0_byteenable               (host_0_lw_bridge_m0_byteenable),        //                               .byteenable
		.lw_bridge_m0_debugaccess              (host_0_lw_bridge_m0_debugaccess),       //                               .debugaccess
		.hps_0_h2f_gp_gp_in                    (host_0_hps_0_h2f_gp_gp_in),             //                   hps_0_h2f_gp.gp_in
		.hps_0_h2f_gp_gp_out                   (host_0_hps_0_h2f_gp_gp_out),            //                               .gp_out
		.hps_0_h2f_cold_reset_reset_n          (host_0_hps_0_h2f_cold_reset_reset_n)    //           hps_0_h2f_cold_reset.reset_n
	);

	soc_system_pcp_0 pcp_0 (
		.clk50_clk                                (clk_50_clk),                          //                             clk50.clk
		.rst_clk50_reset_n                        (reset_reset_n),                       //                         rst_clk50.reset_n
		.clk100_clk                               (clk_100_outclk0_clk),                 //                            clk100.clk
		.rst_clk100_reset_n                       (reset_reset_n),                       //                        rst_clk100.reset_n
		.benchmark_pio_external_connection_export (pcp_0_benchmark_pio_export),          // benchmark_pio_external_connection.export
		.slow_bridge_waitrequest                  (pcp_0_slow_bridge_waitrequest),       //                       slow_bridge.waitrequest
		.slow_bridge_readdata                     (pcp_0_slow_bridge_readdata),          //                                  .readdata
		.slow_bridge_readdatavalid                (pcp_0_slow_bridge_readdatavalid),     //                                  .readdatavalid
		.slow_bridge_burstcount                   (pcp_0_slow_bridge_burstcount),        //                                  .burstcount
		.slow_bridge_writedata                    (pcp_0_slow_bridge_writedata),         //                                  .writedata
		.slow_bridge_address                      (pcp_0_slow_bridge_address),           //                                  .address
		.slow_bridge_write                        (pcp_0_slow_bridge_write),             //                                  .write
		.slow_bridge_read                         (pcp_0_slow_bridge_read),              //                                  .read
		.slow_bridge_byteenable                   (pcp_0_slow_bridge_byteenable),        //                                  .byteenable
		.slow_bridge_debugaccess                  (pcp_0_slow_bridge_debugaccess),       //                                  .debugaccess
		.cpu_bridge_waitrequest                   (pcp_0_cpu_bridge_waitrequest),        //                        cpu_bridge.waitrequest
		.cpu_bridge_readdata                      (pcp_0_cpu_bridge_readdata),           //                                  .readdata
		.cpu_bridge_readdatavalid                 (pcp_0_cpu_bridge_readdatavalid),      //                                  .readdatavalid
		.cpu_bridge_burstcount                    (pcp_0_cpu_bridge_burstcount),         //                                  .burstcount
		.cpu_bridge_writedata                     (pcp_0_cpu_bridge_writedata),          //                                  .writedata
		.cpu_bridge_address                       (pcp_0_cpu_bridge_address),            //                                  .address
		.cpu_bridge_write                         (pcp_0_cpu_bridge_write),              //                                  .write
		.cpu_bridge_read                          (pcp_0_cpu_bridge_read),               //                                  .read
		.cpu_bridge_byteenable                    (pcp_0_cpu_bridge_byteenable),         //                                  .byteenable
		.cpu_bridge_debugaccess                   (pcp_0_cpu_bridge_debugaccess),        //                                  .debugaccess
		.sync_irq_irq                             (pcp_0_sync_irq_irq),                  //                          sync_irq.irq
		.mac_irq_irq                              (pcp_0_mac_irq_irq),                   //                           mac_irq.irq
		.flash_bridge_waitrequest                 (pcp_0_flash_bridge_waitrequest),      //                      flash_bridge.waitrequest
		.flash_bridge_readdata                    (pcp_0_flash_bridge_readdata),         //                                  .readdata
		.flash_bridge_readdatavalid               (pcp_0_flash_bridge_readdatavalid),    //                                  .readdatavalid
		.flash_bridge_burstcount                  (pcp_0_flash_bridge_burstcount),       //                                  .burstcount
		.flash_bridge_writedata                   (pcp_0_flash_bridge_writedata),        //                                  .writedata
		.flash_bridge_address                     (pcp_0_flash_bridge_address),          //                                  .address
		.flash_bridge_write                       (pcp_0_flash_bridge_write),            //                                  .write
		.flash_bridge_read                        (pcp_0_flash_bridge_read),             //                                  .read
		.flash_bridge_byteenable                  (pcp_0_flash_bridge_byteenable),       //                                  .byteenable
		.flash_bridge_debugaccess                 (pcp_0_flash_bridge_debugaccess),      //                                  .debugaccess
		.gp_irq_irq                               (pcp_0_gp_irq_irq),                    //                            gp_irq.irq
		.cpu_resetrequest_resetrequest            (pcp_0_cpu_resetrequest_resetrequest), //                  cpu_resetrequest.resetrequest
		.cpu_resetrequest_resettaken              (pcp_0_cpu_resetrequest_resettaken),   //                                  .resettaken
		.jtag_reset_reset                         (),                                    //                        jtag_reset.reset
		.powerlink_led_export                     (powerlink_led_export)                 //                     powerlink_led.export
	);

	soc_system_mm_interconnect_0 mm_interconnect_0 (
		.clk_100_outclk0_clk                                           (clk_100_outclk0_clk),                                 //                                         clk_100_outclk0.clk
		.clk_50_clk_clk                                                (clk_50_clk),                                          //                                              clk_50_clk.clk
		.host_0_reset_clk50_reset_bridge_in_reset_reset                (rst_controller_reset_out_reset),                      //                host_0_reset_clk50_reset_bridge_in_reset.reset
		.openmac_0_pktBuf_translator_reset_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),                  // openmac_0_pktBuf_translator_reset_reset_bridge_in_reset.reset
		.openmac_0_pktRst_reset_bridge_in_reset_reset                  (rst_controller_001_reset_out_reset),                  //                  openmac_0_pktRst_reset_bridge_in_reset.reset
		.sysid_qsys_reset_reset_bridge_in_reset_reset                  (rst_controller_reset_out_reset),                      //                  sysid_qsys_reset_reset_bridge_in_reset.reset
		.host_0_lw_bridge_m0_address                                   (host_0_lw_bridge_m0_address),                         //                                     host_0_lw_bridge_m0.address
		.host_0_lw_bridge_m0_waitrequest                               (host_0_lw_bridge_m0_waitrequest),                     //                                                        .waitrequest
		.host_0_lw_bridge_m0_burstcount                                (host_0_lw_bridge_m0_burstcount),                      //                                                        .burstcount
		.host_0_lw_bridge_m0_byteenable                                (host_0_lw_bridge_m0_byteenable),                      //                                                        .byteenable
		.host_0_lw_bridge_m0_read                                      (host_0_lw_bridge_m0_read),                            //                                                        .read
		.host_0_lw_bridge_m0_readdata                                  (host_0_lw_bridge_m0_readdata),                        //                                                        .readdata
		.host_0_lw_bridge_m0_readdatavalid                             (host_0_lw_bridge_m0_readdatavalid),                   //                                                        .readdatavalid
		.host_0_lw_bridge_m0_write                                     (host_0_lw_bridge_m0_write),                           //                                                        .write
		.host_0_lw_bridge_m0_writedata                                 (host_0_lw_bridge_m0_writedata),                       //                                                        .writedata
		.host_0_lw_bridge_m0_debugaccess                               (host_0_lw_bridge_m0_debugaccess),                     //                                                        .debugaccess
		.pcp_0_slow_bridge_address                                     (pcp_0_slow_bridge_address),                           //                                       pcp_0_slow_bridge.address
		.pcp_0_slow_bridge_waitrequest                                 (pcp_0_slow_bridge_waitrequest),                       //                                                        .waitrequest
		.pcp_0_slow_bridge_burstcount                                  (pcp_0_slow_bridge_burstcount),                        //                                                        .burstcount
		.pcp_0_slow_bridge_byteenable                                  (pcp_0_slow_bridge_byteenable),                        //                                                        .byteenable
		.pcp_0_slow_bridge_read                                        (pcp_0_slow_bridge_read),                              //                                                        .read
		.pcp_0_slow_bridge_readdata                                    (pcp_0_slow_bridge_readdata),                          //                                                        .readdata
		.pcp_0_slow_bridge_readdatavalid                               (pcp_0_slow_bridge_readdatavalid),                     //                                                        .readdatavalid
		.pcp_0_slow_bridge_write                                       (pcp_0_slow_bridge_write),                             //                                                        .write
		.pcp_0_slow_bridge_writedata                                   (pcp_0_slow_bridge_writedata),                         //                                                        .writedata
		.pcp_0_slow_bridge_debugaccess                                 (pcp_0_slow_bridge_debugaccess),                       //                                                        .debugaccess
		.com_mem_s1_address                                            (mm_interconnect_0_com_mem_s1_address),                //                                              com_mem_s1.address
		.com_mem_s1_write                                              (mm_interconnect_0_com_mem_s1_write),                  //                                                        .write
		.com_mem_s1_readdata                                           (mm_interconnect_0_com_mem_s1_readdata),               //                                                        .readdata
		.com_mem_s1_writedata                                          (mm_interconnect_0_com_mem_s1_writedata),              //                                                        .writedata
		.com_mem_s1_byteenable                                         (mm_interconnect_0_com_mem_s1_byteenable),             //                                                        .byteenable
		.com_mem_s1_chipselect                                         (mm_interconnect_0_com_mem_s1_chipselect),             //                                                        .chipselect
		.com_mem_s1_clken                                              (mm_interconnect_0_com_mem_s1_clken),                  //                                                        .clken
		.com_mem_s2_address                                            (mm_interconnect_0_com_mem_s2_address),                //                                              com_mem_s2.address
		.com_mem_s2_write                                              (mm_interconnect_0_com_mem_s2_write),                  //                                                        .write
		.com_mem_s2_readdata                                           (mm_interconnect_0_com_mem_s2_readdata),               //                                                        .readdata
		.com_mem_s2_writedata                                          (mm_interconnect_0_com_mem_s2_writedata),              //                                                        .writedata
		.com_mem_s2_byteenable                                         (mm_interconnect_0_com_mem_s2_byteenable),             //                                                        .byteenable
		.com_mem_s2_chipselect                                         (mm_interconnect_0_com_mem_s2_chipselect),             //                                                        .chipselect
		.com_mem_s2_clken                                              (mm_interconnect_0_com_mem_s2_clken),                  //                                                        .clken
		.openmac_0_macReg_address                                      (mm_interconnect_0_openmac_0_macreg_address),          //                                        openmac_0_macReg.address
		.openmac_0_macReg_write                                        (mm_interconnect_0_openmac_0_macreg_write),            //                                                        .write
		.openmac_0_macReg_read                                         (mm_interconnect_0_openmac_0_macreg_read),             //                                                        .read
		.openmac_0_macReg_readdata                                     (mm_interconnect_0_openmac_0_macreg_readdata),         //                                                        .readdata
		.openmac_0_macReg_writedata                                    (mm_interconnect_0_openmac_0_macreg_writedata),        //                                                        .writedata
		.openmac_0_macReg_byteenable                                   (mm_interconnect_0_openmac_0_macreg_byteenable),       //                                                        .byteenable
		.openmac_0_macReg_waitrequest                                  (mm_interconnect_0_openmac_0_macreg_waitrequest),      //                                                        .waitrequest
		.openmac_0_macReg_chipselect                                   (mm_interconnect_0_openmac_0_macreg_chipselect),       //                                                        .chipselect
		.openmac_0_macTimer_address                                    (mm_interconnect_0_openmac_0_mactimer_address),        //                                      openmac_0_macTimer.address
		.openmac_0_macTimer_write                                      (mm_interconnect_0_openmac_0_mactimer_write),          //                                                        .write
		.openmac_0_macTimer_read                                       (mm_interconnect_0_openmac_0_mactimer_read),           //                                                        .read
		.openmac_0_macTimer_readdata                                   (mm_interconnect_0_openmac_0_mactimer_readdata),       //                                                        .readdata
		.openmac_0_macTimer_writedata                                  (mm_interconnect_0_openmac_0_mactimer_writedata),      //                                                        .writedata
		.openmac_0_macTimer_byteenable                                 (mm_interconnect_0_openmac_0_mactimer_byteenable),     //                                                        .byteenable
		.openmac_0_macTimer_waitrequest                                (mm_interconnect_0_openmac_0_mactimer_waitrequest),    //                                                        .waitrequest
		.openmac_0_macTimer_chipselect                                 (mm_interconnect_0_openmac_0_mactimer_chipselect),     //                                                        .chipselect
		.openmac_0_pktBuf_address                                      (mm_interconnect_0_openmac_0_pktbuf_address),          //                                        openmac_0_pktBuf.address
		.openmac_0_pktBuf_write                                        (mm_interconnect_0_openmac_0_pktbuf_write),            //                                                        .write
		.openmac_0_pktBuf_read                                         (mm_interconnect_0_openmac_0_pktbuf_read),             //                                                        .read
		.openmac_0_pktBuf_readdata                                     (mm_interconnect_0_openmac_0_pktbuf_readdata),         //                                                        .readdata
		.openmac_0_pktBuf_writedata                                    (mm_interconnect_0_openmac_0_pktbuf_writedata),        //                                                        .writedata
		.openmac_0_pktBuf_byteenable                                   (mm_interconnect_0_openmac_0_pktbuf_byteenable),       //                                                        .byteenable
		.openmac_0_pktBuf_waitrequest                                  (mm_interconnect_0_openmac_0_pktbuf_waitrequest),      //                                                        .waitrequest
		.openmac_0_pktBuf_chipselect                                   (mm_interconnect_0_openmac_0_pktbuf_chipselect),       //                                                        .chipselect
		.sysid_qsys_control_slave_address                              (mm_interconnect_0_sysid_qsys_control_slave_address),  //                                sysid_qsys_control_slave.address
		.sysid_qsys_control_slave_readdata                             (mm_interconnect_0_sysid_qsys_control_slave_readdata)  //                                                        .readdata
	);

	soc_system_mm_interconnect_1 mm_interconnect_1 (
		.clk_100_outclk0_clk                                        (clk_100_outclk0_clk),                              //                                      clk_100_outclk0.clk
		.clk_50_clk_clk                                             (clk_50_clk),                                       //                                           clk_50_clk.clk
		.onchip_memory2_0_reset1_reset_bridge_in_reset_reset        (rst_controller_reset_out_reset),                   //        onchip_memory2_0_reset1_reset_bridge_in_reset.reset
		.openmac_0_dma_translator_reset_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),               // openmac_0_dma_translator_reset_reset_bridge_in_reset.reset
		.openmac_0_dmaRst_reset_bridge_in_reset_reset               (rst_controller_001_reset_out_reset),               //               openmac_0_dmaRst_reset_bridge_in_reset.reset
		.host_0_fpga_mem_address                                    (host_0_fpga_mem_address),                          //                                      host_0_fpga_mem.address
		.host_0_fpga_mem_waitrequest                                (host_0_fpga_mem_waitrequest),                      //                                                     .waitrequest
		.host_0_fpga_mem_burstcount                                 (host_0_fpga_mem_burstcount),                       //                                                     .burstcount
		.host_0_fpga_mem_byteenable                                 (host_0_fpga_mem_byteenable),                       //                                                     .byteenable
		.host_0_fpga_mem_read                                       (host_0_fpga_mem_read),                             //                                                     .read
		.host_0_fpga_mem_readdata                                   (host_0_fpga_mem_readdata),                         //                                                     .readdata
		.host_0_fpga_mem_readdatavalid                              (host_0_fpga_mem_readdatavalid),                    //                                                     .readdatavalid
		.host_0_fpga_mem_write                                      (host_0_fpga_mem_write),                            //                                                     .write
		.host_0_fpga_mem_writedata                                  (host_0_fpga_mem_writedata),                        //                                                     .writedata
		.host_0_fpga_mem_debugaccess                                (host_0_fpga_mem_debugaccess),                      //                                                     .debugaccess
		.openmac_0_dma_address                                      (openmac_0_dma_address),                            //                                        openmac_0_dma.address
		.openmac_0_dma_waitrequest                                  (openmac_0_dma_waitrequest),                        //                                                     .waitrequest
		.openmac_0_dma_burstcount                                   (openmac_0_dma_burstcount),                         //                                                     .burstcount
		.openmac_0_dma_byteenable                                   (openmac_0_dma_byteenable),                         //                                                     .byteenable
		.openmac_0_dma_write                                        (openmac_0_dma_write),                              //                                                     .write
		.openmac_0_dma_writedata                                    (openmac_0_dma_writedata),                          //                                                     .writedata
		.pcp_0_cpu_bridge_address                                   (pcp_0_cpu_bridge_address),                         //                                     pcp_0_cpu_bridge.address
		.pcp_0_cpu_bridge_waitrequest                               (pcp_0_cpu_bridge_waitrequest),                     //                                                     .waitrequest
		.pcp_0_cpu_bridge_burstcount                                (pcp_0_cpu_bridge_burstcount),                      //                                                     .burstcount
		.pcp_0_cpu_bridge_byteenable                                (pcp_0_cpu_bridge_byteenable),                      //                                                     .byteenable
		.pcp_0_cpu_bridge_read                                      (pcp_0_cpu_bridge_read),                            //                                                     .read
		.pcp_0_cpu_bridge_readdata                                  (pcp_0_cpu_bridge_readdata),                        //                                                     .readdata
		.pcp_0_cpu_bridge_readdatavalid                             (pcp_0_cpu_bridge_readdatavalid),                   //                                                     .readdatavalid
		.pcp_0_cpu_bridge_write                                     (pcp_0_cpu_bridge_write),                           //                                                     .write
		.pcp_0_cpu_bridge_writedata                                 (pcp_0_cpu_bridge_writedata),                       //                                                     .writedata
		.pcp_0_cpu_bridge_debugaccess                               (pcp_0_cpu_bridge_debugaccess),                     //                                                     .debugaccess
		.pcp_0_flash_bridge_address                                 (pcp_0_flash_bridge_address),                       //                                   pcp_0_flash_bridge.address
		.pcp_0_flash_bridge_waitrequest                             (pcp_0_flash_bridge_waitrequest),                   //                                                     .waitrequest
		.pcp_0_flash_bridge_burstcount                              (pcp_0_flash_bridge_burstcount),                    //                                                     .burstcount
		.pcp_0_flash_bridge_byteenable                              (pcp_0_flash_bridge_byteenable),                    //                                                     .byteenable
		.pcp_0_flash_bridge_read                                    (pcp_0_flash_bridge_read),                          //                                                     .read
		.pcp_0_flash_bridge_readdata                                (pcp_0_flash_bridge_readdata),                      //                                                     .readdata
		.pcp_0_flash_bridge_readdatavalid                           (pcp_0_flash_bridge_readdatavalid),                 //                                                     .readdatavalid
		.pcp_0_flash_bridge_write                                   (pcp_0_flash_bridge_write),                         //                                                     .write
		.pcp_0_flash_bridge_writedata                               (pcp_0_flash_bridge_writedata),                     //                                                     .writedata
		.pcp_0_flash_bridge_debugaccess                             (pcp_0_flash_bridge_debugaccess),                   //                                                     .debugaccess
		.onchip_memory2_0_s1_address                                (mm_interconnect_1_onchip_memory2_0_s1_address),    //                                  onchip_memory2_0_s1.address
		.onchip_memory2_0_s1_write                                  (mm_interconnect_1_onchip_memory2_0_s1_write),      //                                                     .write
		.onchip_memory2_0_s1_readdata                               (mm_interconnect_1_onchip_memory2_0_s1_readdata),   //                                                     .readdata
		.onchip_memory2_0_s1_writedata                              (mm_interconnect_1_onchip_memory2_0_s1_writedata),  //                                                     .writedata
		.onchip_memory2_0_s1_byteenable                             (mm_interconnect_1_onchip_memory2_0_s1_byteenable), //                                                     .byteenable
		.onchip_memory2_0_s1_chipselect                             (mm_interconnect_1_onchip_memory2_0_s1_chipselect), //                                                     .chipselect
		.onchip_memory2_0_s1_clken                                  (mm_interconnect_1_onchip_memory2_0_s1_clken)       //                                                     .clken
	);

	soc_system_irq_mapper irq_mapper (
		.clk           (clk_50_clk),               //       clk.clk
		.reset         (),                         // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq), // receiver0.irq
		.sender_irq    (host_0_hostif_irq_i_irq)   //    sender.irq
	);

	soc_system_irq_mapper irq_mapper_001 (
		.clk           (clk_50_clk),                     //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_001_receiver0_irq),   // receiver0.irq
		.sender_irq    (pcp_0_sync_irq_irq)              //    sender.irq
	);

	soc_system_irq_mapper irq_mapper_002 (
		.clk           (clk_50_clk),                     //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_002_receiver0_irq),   // receiver0.irq
		.sender_irq    (pcp_0_mac_irq_irq)               //    sender.irq
	);

	soc_system_irq_mapper_003 irq_mapper_003 (
		.clk        (clk_50_clk),                     //       clk.clk
		.reset      (rst_controller_reset_out_reset), // clk_reset.reset
		.sender_irq (pcp_0_gp_irq_irq)                //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (clk_50_clk),                         //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (clk_100_outclk0_clk),                //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
