// mn_soc_host_de10_nano_soc.v

// Generated using ACDS version 14.0 200 at 2018.01.25.20:11:59

`timescale 1 ps / 1 ps
module mn_soc_host_de10_nano_soc (
		output wire [14:0] memory_mem_a,                                           //                                 memory.mem_a
		output wire [2:0]  memory_mem_ba,                                          //                                       .mem_ba
		output wire        memory_mem_ck,                                          //                                       .mem_ck
		output wire        memory_mem_ck_n,                                        //                                       .mem_ck_n
		output wire        memory_mem_cke,                                         //                                       .mem_cke
		output wire        memory_mem_cs_n,                                        //                                       .mem_cs_n
		output wire        memory_mem_ras_n,                                       //                                       .mem_ras_n
		output wire        memory_mem_cas_n,                                       //                                       .mem_cas_n
		output wire        memory_mem_we_n,                                        //                                       .mem_we_n
		output wire        memory_mem_reset_n,                                     //                                       .mem_reset_n
		inout  wire [31:0] memory_mem_dq,                                          //                                       .mem_dq
		inout  wire [3:0]  memory_mem_dqs,                                         //                                       .mem_dqs
		inout  wire [3:0]  memory_mem_dqs_n,                                       //                                       .mem_dqs_n
		output wire        memory_mem_odt,                                         //                                       .mem_odt
		output wire [3:0]  memory_mem_dm,                                          //                                       .mem_dm
		input  wire        memory_oct_rzqin,                                       //                                       .oct_rzqin
		input  wire        clk50_clk,                                              //                                  clk50.clk
		input  wire        reset_clk50_reset_n,                                    //                            reset_clk50.reset_n
		inout  wire        hps_0_hps_io_hps_io_sdio_inst_CMD,                      //                           hps_0_hps_io.hps_io_sdio_inst_CMD
		inout  wire        hps_0_hps_io_hps_io_sdio_inst_D0,                       //                                       .hps_io_sdio_inst_D0
		inout  wire        hps_0_hps_io_hps_io_sdio_inst_D1,                       //                                       .hps_io_sdio_inst_D1
		output wire        hps_0_hps_io_hps_io_sdio_inst_CLK,                      //                                       .hps_io_sdio_inst_CLK
		inout  wire        hps_0_hps_io_hps_io_sdio_inst_D2,                       //                                       .hps_io_sdio_inst_D2
		inout  wire        hps_0_hps_io_hps_io_sdio_inst_D3,                       //                                       .hps_io_sdio_inst_D3
		inout  wire        hps_0_hps_io_hps_io_usb1_inst_D0,                       //                                       .hps_io_usb1_inst_D0
		inout  wire        hps_0_hps_io_hps_io_usb1_inst_D1,                       //                                       .hps_io_usb1_inst_D1
		inout  wire        hps_0_hps_io_hps_io_usb1_inst_D2,                       //                                       .hps_io_usb1_inst_D2
		inout  wire        hps_0_hps_io_hps_io_usb1_inst_D3,                       //                                       .hps_io_usb1_inst_D3
		inout  wire        hps_0_hps_io_hps_io_usb1_inst_D4,                       //                                       .hps_io_usb1_inst_D4
		inout  wire        hps_0_hps_io_hps_io_usb1_inst_D5,                       //                                       .hps_io_usb1_inst_D5
		inout  wire        hps_0_hps_io_hps_io_usb1_inst_D6,                       //                                       .hps_io_usb1_inst_D6
		inout  wire        hps_0_hps_io_hps_io_usb1_inst_D7,                       //                                       .hps_io_usb1_inst_D7
		input  wire        hps_0_hps_io_hps_io_usb1_inst_CLK,                      //                                       .hps_io_usb1_inst_CLK
		output wire        hps_0_hps_io_hps_io_usb1_inst_STP,                      //                                       .hps_io_usb1_inst_STP
		input  wire        hps_0_hps_io_hps_io_usb1_inst_DIR,                      //                                       .hps_io_usb1_inst_DIR
		input  wire        hps_0_hps_io_hps_io_usb1_inst_NXT,                      //                                       .hps_io_usb1_inst_NXT
		output wire        hps_0_hps_io_hps_io_spim1_inst_CLK,                     //                                       .hps_io_spim1_inst_CLK
		output wire        hps_0_hps_io_hps_io_spim1_inst_MOSI,                    //                                       .hps_io_spim1_inst_MOSI
		input  wire        hps_0_hps_io_hps_io_spim1_inst_MISO,                    //                                       .hps_io_spim1_inst_MISO
		output wire        hps_0_hps_io_hps_io_spim1_inst_SS0,                     //                                       .hps_io_spim1_inst_SS0
		input  wire        hps_0_hps_io_hps_io_uart0_inst_RX,                      //                                       .hps_io_uart0_inst_RX
		output wire        hps_0_hps_io_hps_io_uart0_inst_TX,                      //                                       .hps_io_uart0_inst_TX
		inout  wire        hps_0_hps_io_hps_io_i2c0_inst_SDA,                      //                                       .hps_io_i2c0_inst_SDA
		inout  wire        hps_0_hps_io_hps_io_i2c0_inst_SCL,                      //                                       .hps_io_i2c0_inst_SCL
		inout  wire        hps_0_hps_io_hps_io_i2c1_inst_SDA,                      //                                       .hps_io_i2c1_inst_SDA
		inout  wire        hps_0_hps_io_hps_io_i2c1_inst_SCL,                      //                                       .hps_io_i2c1_inst_SCL
		inout  wire        hps_0_hps_io_hps_io_gpio_inst_GPIO09,                   //                                       .hps_io_gpio_inst_GPIO09
		inout  wire        hps_0_hps_io_hps_io_gpio_inst_GPIO35,                   //                                       .hps_io_gpio_inst_GPIO35
		inout  wire        hps_0_hps_io_hps_io_gpio_inst_GPIO40,                   //                                       .hps_io_gpio_inst_GPIO40
		inout  wire        hps_0_hps_io_hps_io_gpio_inst_GPIO53,                   //                                       .hps_io_gpio_inst_GPIO53
		inout  wire        hps_0_hps_io_hps_io_gpio_inst_GPIO54,                   //                                       .hps_io_gpio_inst_GPIO54
		inout  wire        hps_0_hps_io_hps_io_gpio_inst_GPIO61,                   //                                       .hps_io_gpio_inst_GPIO61
		inout  wire        hps_0_hps_io_hps_io_gpio_inst_LOANIO20,                 //                                       .hps_io_gpio_inst_LOANIO20
		inout  wire        hps_0_hps_io_hps_io_gpio_inst_LOANIO21,                 //                                       .hps_io_gpio_inst_LOANIO21
		input  wire [3:0]  dipsw_pio_external_connection_export,                   //          dipsw_pio_external_connection.export
		input  wire [1:0]  button_pio_external_connection_export,                  //         button_pio_external_connection.export
		input  wire        hps_0_f2h_cold_reset_req_reset_n,                       //               hps_0_f2h_cold_reset_req.reset_n
		input  wire        hps_0_f2h_debug_reset_req_reset_n,                      //              hps_0_f2h_debug_reset_req.reset_n
		input  wire        hps_0_f2h_warm_reset_req_reset_n,                       //               hps_0_f2h_warm_reset_req.reset_n
		input  wire        clk100_clk,                                             //                                 clk100.clk
		input  wire        fpga_mem_waitrequest,                                   //                               fpga_mem.waitrequest
		input  wire [31:0] fpga_mem_readdata,                                      //                                       .readdata
		input  wire        fpga_mem_readdatavalid,                                 //                                       .readdatavalid
		output wire [0:0]  fpga_mem_burstcount,                                    //                                       .burstcount
		output wire [31:0] fpga_mem_writedata,                                     //                                       .writedata
		output wire [26:0] fpga_mem_address,                                       //                                       .address
		output wire        fpga_mem_write,                                         //                                       .write
		output wire        fpga_mem_read,                                          //                                       .read
		output wire [3:0]  fpga_mem_byteenable,                                    //                                       .byteenable
		output wire        fpga_mem_debugaccess,                                   //                                       .debugaccess
		input  wire        reset_clk100_reset_n,                                   //                           reset_clk100.reset_n
		input  wire [0:0]  hostif_irq_i_irq,                                       //                           hostif_irq_i.irq
		input  wire        lw_bridge_m0_waitrequest,                               //                           lw_bridge_m0.waitrequest
		input  wire [31:0] lw_bridge_m0_readdata,                                  //                                       .readdata
		input  wire        lw_bridge_m0_readdatavalid,                             //                                       .readdatavalid
		output wire [0:0]  lw_bridge_m0_burstcount,                                //                                       .burstcount
		output wire [31:0] lw_bridge_m0_writedata,                                 //                                       .writedata
		output wire [17:0] lw_bridge_m0_address,                                   //                                       .address
		output wire        lw_bridge_m0_write,                                     //                                       .write
		output wire        lw_bridge_m0_read,                                      //                                       .read
		output wire [3:0]  lw_bridge_m0_byteenable,                                //                                       .byteenable
		output wire        lw_bridge_m0_debugaccess,                               //                                       .debugaccess
		input  wire [31:0] hps_0_h2f_gp_gp_in,                                     //                           hps_0_h2f_gp.gp_in
		output wire [31:0] hps_0_h2f_gp_gp_out,                                    //                                       .gp_out
		output wire        hps_0_h2f_cold_reset_reset_n,                           //                   hps_0_h2f_cold_reset.reset_n
		output wire [66:0] hps_0_h2f_loan_io_in,                                   //                      hps_0_h2f_loan_io.in
		input  wire [66:0] hps_0_h2f_loan_io_out,                                  //                                       .out
		input  wire [66:0] hps_0_h2f_loan_io_oe,                                   //                                       .oe
		output wire        hps_0_emac1_md_clk_clk,                                 //                     hps_0_emac1_md_clk.clk
		input  wire        hps_emac_interface_splitter_0_hps_gmii_phy_tx_clk_i,    // hps_emac_interface_splitter_0_hps_gmii.phy_tx_clk_i
		input  wire        hps_emac_interface_splitter_0_hps_gmii_phy_rx_clk_i,    //                                       .phy_rx_clk_i
		input  wire        hps_emac_interface_splitter_0_hps_gmii_phy_rxdv_i,      //                                       .phy_rxdv_i
		input  wire        hps_emac_interface_splitter_0_hps_gmii_phy_rxer_i,      //                                       .phy_rxer_i
		input  wire [7:0]  hps_emac_interface_splitter_0_hps_gmii_phy_rxd_i,       //                                       .phy_rxd_i
		input  wire        hps_emac_interface_splitter_0_hps_gmii_phy_col_i,       //                                       .phy_col_i
		input  wire        hps_emac_interface_splitter_0_hps_gmii_phy_crs_i,       //                                       .phy_crs_i
		output wire        hps_emac_interface_splitter_0_hps_gmii_phy_tx_clk_o,    //                                       .phy_tx_clk_o
		output wire        hps_emac_interface_splitter_0_hps_gmii_rst_tx_n,        //                                       .rst_tx_n
		output wire        hps_emac_interface_splitter_0_hps_gmii_rst_rx_n,        //                                       .rst_rx_n
		output wire [7:0]  hps_emac_interface_splitter_0_hps_gmii_phy_txd_o,       //                                       .phy_txd_o
		output wire        hps_emac_interface_splitter_0_hps_gmii_phy_txen_o,      //                                       .phy_txen_o
		output wire        hps_emac_interface_splitter_0_hps_gmii_phy_txer_o,      //                                       .phy_txer_o
		output wire [1:0]  hps_emac_interface_splitter_0_hps_gmii_phy_mac_speed_o, //                                       .phy_mac_speed_o
		input  wire        hps_emac_interface_splitter_0_ptp_ptp_aux_ts_trig_i,    //      hps_emac_interface_splitter_0_ptp.ptp_aux_ts_trig_i
		output wire        hps_emac_interface_splitter_0_ptp_ptp_pps_o,            //                                       .ptp_pps_o
		input  wire        hps_emac_interface_splitter_0_mdio_gmii_mdi_i,          //     hps_emac_interface_splitter_0_mdio.gmii_mdi_i
		output wire        hps_emac_interface_splitter_0_mdio_gmii_mdo_o,          //                                       .gmii_mdo_o
		output wire        hps_emac_interface_splitter_0_mdio_gmii_mdo_o_e         //                                       .gmii_mdo_o_e
	);

	wire         hps_emac_interface_splitter_0_emac_phy_crs_i;                // hps_emac_interface_splitter_0:phy_crs_i -> hps_0:emac1_phy_crs_i
	wire   [7:0] hps_emac_interface_splitter_0_emac_phy_rxd_i;                // hps_emac_interface_splitter_0:phy_rxd_i -> hps_0:emac1_phy_rxd_i
	wire         hps_emac_interface_splitter_0_emac_gmii_mdi_i;               // hps_emac_interface_splitter_0:mdi_i -> hps_0:emac1_gmii_mdi_i
	wire         hps_emac_interface_splitter_0_emac_phy_col_i;                // hps_emac_interface_splitter_0:phy_col_i -> hps_0:emac1_phy_col_i
	wire         hps_0_emac1_gmii_mdo_o;                                      // hps_0:emac1_gmii_mdo_o -> hps_emac_interface_splitter_0:mdo_o
	wire         hps_0_emac1_ptp_pps_o;                                       // hps_0:emac1_ptp_pps_o -> hps_emac_interface_splitter_0:ptp_pps_o
	wire   [7:0] hps_0_emac1_phy_txd_o;                                       // hps_0:emac1_phy_txd_o -> hps_emac_interface_splitter_0:phy_txd_o
	wire         hps_0_emac1_phy_txen_o;                                      // hps_0:emac1_phy_txen_o -> hps_emac_interface_splitter_0:phy_txen_o
	wire         hps_emac_interface_splitter_0_emac_phy_rxer_i;               // hps_emac_interface_splitter_0:phy_rxer_i -> hps_0:emac1_phy_rxer_i
	wire         hps_0_emac1_phy_txer_o;                                      // hps_0:emac1_phy_txer_o -> hps_emac_interface_splitter_0:phy_txer_o
	wire         hps_0_emac1_gmii_mdo_o_e;                                    // hps_0:emac1_gmii_mdo_o_e -> hps_emac_interface_splitter_0:mdo_o_e
	wire         hps_emac_interface_splitter_0_emac_ptp_aux_ts_trig_i;        // hps_emac_interface_splitter_0:ptp_aux_ts_trig_i -> hps_0:emac1_ptp_aux_ts_trig_i
	wire         hps_emac_interface_splitter_0_emac_phy_rxdv_i;               // hps_emac_interface_splitter_0:phy_rxdv_i -> hps_0:emac1_phy_rxdv_i
	wire         hps_0_emac1_gtx_clk_clk;                                     // hps_0:emac1_phy_txclk_o -> [hps_emac_interface_splitter_0:phy_txclk_o, rst_controller_003:clk]
	wire         hps_emac_interface_splitter_0_emac_tx_clk_in_clk;            // hps_emac_interface_splitter_0:clk_tx_i -> hps_0:emac1_clk_tx_i
	wire         hps_emac_interface_splitter_0_emac_rx_clk_in_clk;            // hps_emac_interface_splitter_0:clk_rx_i -> hps_0:emac1_clk_rx_i
	wire         hps_0_emac1_rx_reset_reset;                                  // hps_0:emac1_rst_clk_rx_n_o -> hps_emac_interface_splitter_0:rst_rx_n_o
	wire         hps_0_h2f_lw_axi_master_awvalid;                             // hps_0:h2f_lw_AWVALID -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awvalid
	wire   [2:0] hps_0_h2f_lw_axi_master_arsize;                              // hps_0:h2f_lw_ARSIZE -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arsize
	wire   [1:0] hps_0_h2f_lw_axi_master_arlock;                              // hps_0:h2f_lw_ARLOCK -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arlock
	wire   [3:0] hps_0_h2f_lw_axi_master_awcache;                             // hps_0:h2f_lw_AWCACHE -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awcache
	wire         hps_0_h2f_lw_axi_master_arready;                             // mm_interconnect_0:hps_0_h2f_lw_axi_master_arready -> hps_0:h2f_lw_ARREADY
	wire  [11:0] hps_0_h2f_lw_axi_master_arid;                                // hps_0:h2f_lw_ARID -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arid
	wire         hps_0_h2f_lw_axi_master_rready;                              // hps_0:h2f_lw_RREADY -> mm_interconnect_0:hps_0_h2f_lw_axi_master_rready
	wire         hps_0_h2f_lw_axi_master_bready;                              // hps_0:h2f_lw_BREADY -> mm_interconnect_0:hps_0_h2f_lw_axi_master_bready
	wire   [2:0] hps_0_h2f_lw_axi_master_awsize;                              // hps_0:h2f_lw_AWSIZE -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awsize
	wire   [2:0] hps_0_h2f_lw_axi_master_awprot;                              // hps_0:h2f_lw_AWPROT -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awprot
	wire         hps_0_h2f_lw_axi_master_arvalid;                             // hps_0:h2f_lw_ARVALID -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arvalid
	wire   [2:0] hps_0_h2f_lw_axi_master_arprot;                              // hps_0:h2f_lw_ARPROT -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arprot
	wire  [11:0] hps_0_h2f_lw_axi_master_bid;                                 // mm_interconnect_0:hps_0_h2f_lw_axi_master_bid -> hps_0:h2f_lw_BID
	wire   [3:0] hps_0_h2f_lw_axi_master_arlen;                               // hps_0:h2f_lw_ARLEN -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arlen
	wire         hps_0_h2f_lw_axi_master_awready;                             // mm_interconnect_0:hps_0_h2f_lw_axi_master_awready -> hps_0:h2f_lw_AWREADY
	wire  [11:0] hps_0_h2f_lw_axi_master_awid;                                // hps_0:h2f_lw_AWID -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awid
	wire         hps_0_h2f_lw_axi_master_bvalid;                              // mm_interconnect_0:hps_0_h2f_lw_axi_master_bvalid -> hps_0:h2f_lw_BVALID
	wire  [11:0] hps_0_h2f_lw_axi_master_wid;                                 // hps_0:h2f_lw_WID -> mm_interconnect_0:hps_0_h2f_lw_axi_master_wid
	wire   [1:0] hps_0_h2f_lw_axi_master_awlock;                              // hps_0:h2f_lw_AWLOCK -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awlock
	wire   [1:0] hps_0_h2f_lw_axi_master_awburst;                             // hps_0:h2f_lw_AWBURST -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awburst
	wire   [1:0] hps_0_h2f_lw_axi_master_bresp;                               // mm_interconnect_0:hps_0_h2f_lw_axi_master_bresp -> hps_0:h2f_lw_BRESP
	wire   [3:0] hps_0_h2f_lw_axi_master_wstrb;                               // hps_0:h2f_lw_WSTRB -> mm_interconnect_0:hps_0_h2f_lw_axi_master_wstrb
	wire         hps_0_h2f_lw_axi_master_rvalid;                              // mm_interconnect_0:hps_0_h2f_lw_axi_master_rvalid -> hps_0:h2f_lw_RVALID
	wire  [31:0] hps_0_h2f_lw_axi_master_wdata;                               // hps_0:h2f_lw_WDATA -> mm_interconnect_0:hps_0_h2f_lw_axi_master_wdata
	wire         hps_0_h2f_lw_axi_master_wready;                              // mm_interconnect_0:hps_0_h2f_lw_axi_master_wready -> hps_0:h2f_lw_WREADY
	wire   [1:0] hps_0_h2f_lw_axi_master_arburst;                             // hps_0:h2f_lw_ARBURST -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arburst
	wire  [31:0] hps_0_h2f_lw_axi_master_rdata;                               // mm_interconnect_0:hps_0_h2f_lw_axi_master_rdata -> hps_0:h2f_lw_RDATA
	wire  [20:0] hps_0_h2f_lw_axi_master_araddr;                              // hps_0:h2f_lw_ARADDR -> mm_interconnect_0:hps_0_h2f_lw_axi_master_araddr
	wire   [3:0] hps_0_h2f_lw_axi_master_arcache;                             // hps_0:h2f_lw_ARCACHE -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arcache
	wire   [3:0] hps_0_h2f_lw_axi_master_awlen;                               // hps_0:h2f_lw_AWLEN -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awlen
	wire  [20:0] hps_0_h2f_lw_axi_master_awaddr;                              // hps_0:h2f_lw_AWADDR -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awaddr
	wire  [11:0] hps_0_h2f_lw_axi_master_rid;                                 // mm_interconnect_0:hps_0_h2f_lw_axi_master_rid -> hps_0:h2f_lw_RID
	wire         hps_0_h2f_lw_axi_master_wvalid;                              // hps_0:h2f_lw_WVALID -> mm_interconnect_0:hps_0_h2f_lw_axi_master_wvalid
	wire   [1:0] hps_0_h2f_lw_axi_master_rresp;                               // mm_interconnect_0:hps_0_h2f_lw_axi_master_rresp -> hps_0:h2f_lw_RRESP
	wire         hps_0_h2f_lw_axi_master_wlast;                               // hps_0:h2f_lw_WLAST -> mm_interconnect_0:hps_0_h2f_lw_axi_master_wlast
	wire         hps_0_h2f_lw_axi_master_rlast;                               // mm_interconnect_0:hps_0_h2f_lw_axi_master_rlast -> hps_0:h2f_lw_RLAST
	wire  [31:0] mm_interconnect_0_dipsw_pio_s1_writedata;                    // mm_interconnect_0:dipsw_pio_s1_writedata -> dipsw_pio:writedata
	wire   [1:0] mm_interconnect_0_dipsw_pio_s1_address;                      // mm_interconnect_0:dipsw_pio_s1_address -> dipsw_pio:address
	wire         mm_interconnect_0_dipsw_pio_s1_chipselect;                   // mm_interconnect_0:dipsw_pio_s1_chipselect -> dipsw_pio:chipselect
	wire         mm_interconnect_0_dipsw_pio_s1_write;                        // mm_interconnect_0:dipsw_pio_s1_write -> dipsw_pio:write_n
	wire  [31:0] mm_interconnect_0_dipsw_pio_s1_readdata;                     // dipsw_pio:readdata -> mm_interconnect_0:dipsw_pio_s1_readdata
	wire  [31:0] mm_interconnect_0_button_pio_s1_writedata;                   // mm_interconnect_0:button_pio_s1_writedata -> button_pio:writedata
	wire   [1:0] mm_interconnect_0_button_pio_s1_address;                     // mm_interconnect_0:button_pio_s1_address -> button_pio:address
	wire         mm_interconnect_0_button_pio_s1_chipselect;                  // mm_interconnect_0:button_pio_s1_chipselect -> button_pio:chipselect
	wire         mm_interconnect_0_button_pio_s1_write;                       // mm_interconnect_0:button_pio_s1_write -> button_pio:write_n
	wire  [31:0] mm_interconnect_0_button_pio_s1_readdata;                    // button_pio:readdata -> mm_interconnect_0:button_pio_s1_readdata
	wire         mm_interconnect_0_lw_bridge_s0_waitrequest;                  // lw_bridge:s0_waitrequest -> mm_interconnect_0:lw_bridge_s0_waitrequest
	wire   [0:0] mm_interconnect_0_lw_bridge_s0_burstcount;                   // mm_interconnect_0:lw_bridge_s0_burstcount -> lw_bridge:s0_burstcount
	wire  [31:0] mm_interconnect_0_lw_bridge_s0_writedata;                    // mm_interconnect_0:lw_bridge_s0_writedata -> lw_bridge:s0_writedata
	wire  [17:0] mm_interconnect_0_lw_bridge_s0_address;                      // mm_interconnect_0:lw_bridge_s0_address -> lw_bridge:s0_address
	wire         mm_interconnect_0_lw_bridge_s0_write;                        // mm_interconnect_0:lw_bridge_s0_write -> lw_bridge:s0_write
	wire         mm_interconnect_0_lw_bridge_s0_read;                         // mm_interconnect_0:lw_bridge_s0_read -> lw_bridge:s0_read
	wire  [31:0] mm_interconnect_0_lw_bridge_s0_readdata;                     // lw_bridge:s0_readdata -> mm_interconnect_0:lw_bridge_s0_readdata
	wire         mm_interconnect_0_lw_bridge_s0_debugaccess;                  // mm_interconnect_0:lw_bridge_s0_debugaccess -> lw_bridge:s0_debugaccess
	wire         mm_interconnect_0_lw_bridge_s0_readdatavalid;                // lw_bridge:s0_readdatavalid -> mm_interconnect_0:lw_bridge_s0_readdatavalid
	wire   [3:0] mm_interconnect_0_lw_bridge_s0_byteenable;                   // mm_interconnect_0:lw_bridge_s0_byteenable -> lw_bridge:s0_byteenable
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest; // jtag_uart_0:av_waitrequest -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_waitrequest
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata;   // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_writedata -> jtag_uart_0:av_writedata
	wire   [0:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address;     // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_address -> jtag_uart_0:av_address
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect;  // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_chipselect -> jtag_uart_0:av_chipselect
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write;       // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_write -> jtag_uart_0:av_write_n
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read;        // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_read -> jtag_uart_0:av_read_n
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata;    // jtag_uart_0:av_readdata -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_readdata
	wire  [15:0] mm_interconnect_0_timer_0_s1_writedata;                      // mm_interconnect_0:timer_0_s1_writedata -> timer_0:writedata
	wire   [2:0] mm_interconnect_0_timer_0_s1_address;                        // mm_interconnect_0:timer_0_s1_address -> timer_0:address
	wire         mm_interconnect_0_timer_0_s1_chipselect;                     // mm_interconnect_0:timer_0_s1_chipselect -> timer_0:chipselect
	wire         mm_interconnect_0_timer_0_s1_write;                          // mm_interconnect_0:timer_0_s1_write -> timer_0:write_n
	wire  [15:0] mm_interconnect_0_timer_0_s1_readdata;                       // timer_0:readdata -> mm_interconnect_0:timer_0_s1_readdata
	wire         hps_0_h2f_axi_master_awvalid;                                // hps_0:h2f_AWVALID -> mm_interconnect_1:hps_0_h2f_axi_master_awvalid
	wire   [2:0] hps_0_h2f_axi_master_arsize;                                 // hps_0:h2f_ARSIZE -> mm_interconnect_1:hps_0_h2f_axi_master_arsize
	wire   [1:0] hps_0_h2f_axi_master_arlock;                                 // hps_0:h2f_ARLOCK -> mm_interconnect_1:hps_0_h2f_axi_master_arlock
	wire   [3:0] hps_0_h2f_axi_master_awcache;                                // hps_0:h2f_AWCACHE -> mm_interconnect_1:hps_0_h2f_axi_master_awcache
	wire         hps_0_h2f_axi_master_arready;                                // mm_interconnect_1:hps_0_h2f_axi_master_arready -> hps_0:h2f_ARREADY
	wire  [11:0] hps_0_h2f_axi_master_arid;                                   // hps_0:h2f_ARID -> mm_interconnect_1:hps_0_h2f_axi_master_arid
	wire         hps_0_h2f_axi_master_rready;                                 // hps_0:h2f_RREADY -> mm_interconnect_1:hps_0_h2f_axi_master_rready
	wire         hps_0_h2f_axi_master_bready;                                 // hps_0:h2f_BREADY -> mm_interconnect_1:hps_0_h2f_axi_master_bready
	wire   [2:0] hps_0_h2f_axi_master_awsize;                                 // hps_0:h2f_AWSIZE -> mm_interconnect_1:hps_0_h2f_axi_master_awsize
	wire   [2:0] hps_0_h2f_axi_master_awprot;                                 // hps_0:h2f_AWPROT -> mm_interconnect_1:hps_0_h2f_axi_master_awprot
	wire         hps_0_h2f_axi_master_arvalid;                                // hps_0:h2f_ARVALID -> mm_interconnect_1:hps_0_h2f_axi_master_arvalid
	wire   [2:0] hps_0_h2f_axi_master_arprot;                                 // hps_0:h2f_ARPROT -> mm_interconnect_1:hps_0_h2f_axi_master_arprot
	wire  [11:0] hps_0_h2f_axi_master_bid;                                    // mm_interconnect_1:hps_0_h2f_axi_master_bid -> hps_0:h2f_BID
	wire   [3:0] hps_0_h2f_axi_master_arlen;                                  // hps_0:h2f_ARLEN -> mm_interconnect_1:hps_0_h2f_axi_master_arlen
	wire         hps_0_h2f_axi_master_awready;                                // mm_interconnect_1:hps_0_h2f_axi_master_awready -> hps_0:h2f_AWREADY
	wire  [11:0] hps_0_h2f_axi_master_awid;                                   // hps_0:h2f_AWID -> mm_interconnect_1:hps_0_h2f_axi_master_awid
	wire         hps_0_h2f_axi_master_bvalid;                                 // mm_interconnect_1:hps_0_h2f_axi_master_bvalid -> hps_0:h2f_BVALID
	wire  [11:0] hps_0_h2f_axi_master_wid;                                    // hps_0:h2f_WID -> mm_interconnect_1:hps_0_h2f_axi_master_wid
	wire   [1:0] hps_0_h2f_axi_master_awlock;                                 // hps_0:h2f_AWLOCK -> mm_interconnect_1:hps_0_h2f_axi_master_awlock
	wire   [1:0] hps_0_h2f_axi_master_awburst;                                // hps_0:h2f_AWBURST -> mm_interconnect_1:hps_0_h2f_axi_master_awburst
	wire   [1:0] hps_0_h2f_axi_master_bresp;                                  // mm_interconnect_1:hps_0_h2f_axi_master_bresp -> hps_0:h2f_BRESP
	wire   [3:0] hps_0_h2f_axi_master_wstrb;                                  // hps_0:h2f_WSTRB -> mm_interconnect_1:hps_0_h2f_axi_master_wstrb
	wire         hps_0_h2f_axi_master_rvalid;                                 // mm_interconnect_1:hps_0_h2f_axi_master_rvalid -> hps_0:h2f_RVALID
	wire  [31:0] hps_0_h2f_axi_master_wdata;                                  // hps_0:h2f_WDATA -> mm_interconnect_1:hps_0_h2f_axi_master_wdata
	wire         hps_0_h2f_axi_master_wready;                                 // mm_interconnect_1:hps_0_h2f_axi_master_wready -> hps_0:h2f_WREADY
	wire   [1:0] hps_0_h2f_axi_master_arburst;                                // hps_0:h2f_ARBURST -> mm_interconnect_1:hps_0_h2f_axi_master_arburst
	wire  [31:0] hps_0_h2f_axi_master_rdata;                                  // mm_interconnect_1:hps_0_h2f_axi_master_rdata -> hps_0:h2f_RDATA
	wire  [29:0] hps_0_h2f_axi_master_araddr;                                 // hps_0:h2f_ARADDR -> mm_interconnect_1:hps_0_h2f_axi_master_araddr
	wire   [3:0] hps_0_h2f_axi_master_arcache;                                // hps_0:h2f_ARCACHE -> mm_interconnect_1:hps_0_h2f_axi_master_arcache
	wire   [3:0] hps_0_h2f_axi_master_awlen;                                  // hps_0:h2f_AWLEN -> mm_interconnect_1:hps_0_h2f_axi_master_awlen
	wire  [29:0] hps_0_h2f_axi_master_awaddr;                                 // hps_0:h2f_AWADDR -> mm_interconnect_1:hps_0_h2f_axi_master_awaddr
	wire  [11:0] hps_0_h2f_axi_master_rid;                                    // mm_interconnect_1:hps_0_h2f_axi_master_rid -> hps_0:h2f_RID
	wire         hps_0_h2f_axi_master_wvalid;                                 // hps_0:h2f_WVALID -> mm_interconnect_1:hps_0_h2f_axi_master_wvalid
	wire   [1:0] hps_0_h2f_axi_master_rresp;                                  // mm_interconnect_1:hps_0_h2f_axi_master_rresp -> hps_0:h2f_RRESP
	wire         hps_0_h2f_axi_master_wlast;                                  // hps_0:h2f_WLAST -> mm_interconnect_1:hps_0_h2f_axi_master_wlast
	wire         hps_0_h2f_axi_master_rlast;                                  // mm_interconnect_1:hps_0_h2f_axi_master_rlast -> hps_0:h2f_RLAST
	wire         mm_interconnect_1_fpga_mem_s0_waitrequest;                   // fpga_mem:s0_waitrequest -> mm_interconnect_1:fpga_mem_s0_waitrequest
	wire   [0:0] mm_interconnect_1_fpga_mem_s0_burstcount;                    // mm_interconnect_1:fpga_mem_s0_burstcount -> fpga_mem:s0_burstcount
	wire  [31:0] mm_interconnect_1_fpga_mem_s0_writedata;                     // mm_interconnect_1:fpga_mem_s0_writedata -> fpga_mem:s0_writedata
	wire  [26:0] mm_interconnect_1_fpga_mem_s0_address;                       // mm_interconnect_1:fpga_mem_s0_address -> fpga_mem:s0_address
	wire         mm_interconnect_1_fpga_mem_s0_write;                         // mm_interconnect_1:fpga_mem_s0_write -> fpga_mem:s0_write
	wire         mm_interconnect_1_fpga_mem_s0_read;                          // mm_interconnect_1:fpga_mem_s0_read -> fpga_mem:s0_read
	wire  [31:0] mm_interconnect_1_fpga_mem_s0_readdata;                      // fpga_mem:s0_readdata -> mm_interconnect_1:fpga_mem_s0_readdata
	wire         mm_interconnect_1_fpga_mem_s0_debugaccess;                   // mm_interconnect_1:fpga_mem_s0_debugaccess -> fpga_mem:s0_debugaccess
	wire         mm_interconnect_1_fpga_mem_s0_readdatavalid;                 // fpga_mem:s0_readdatavalid -> mm_interconnect_1:fpga_mem_s0_readdatavalid
	wire   [3:0] mm_interconnect_1_fpga_mem_s0_byteenable;                    // mm_interconnect_1:fpga_mem_s0_byteenable -> fpga_mem:s0_byteenable
	wire         irq_mapper_receiver0_irq;                                    // hostif_irq:sender0_irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                    // jtag_uart_0:av_irq -> irq_mapper:receiver1_irq
	wire         irq_mapper_receiver2_irq;                                    // timer_0:irq -> irq_mapper:receiver2_irq
	wire  [31:0] hps_0_f2h_irq0_irq;                                          // irq_mapper:sender_irq -> hps_0:f2h_irq_p0
	wire  [31:0] hps_0_f2h_irq1_irq;                                          // irq_mapper_001:sender_irq -> hps_0:f2h_irq_p1
	wire         rst_controller_reset_out_reset;                              // rst_controller:reset_out -> [button_pio:reset_n, dipsw_pio:reset_n, hps_emac_interface_splitter_0:rst_n, jtag_uart_0:rst_n, mm_interconnect_0:dipsw_pio_reset_reset_bridge_in_reset_reset]
	wire         rst_controller_001_reset_out_reset;                          // rst_controller_001:reset_out -> [fpga_mem:reset, mm_interconnect_1:fpga_mem_reset_reset_bridge_in_reset_reset]
	wire         rst_controller_002_reset_out_reset;                          // rst_controller_002:reset_out -> [hostif_irq:reset, lw_bridge:reset, mm_interconnect_0:lw_bridge_reset_reset_bridge_in_reset_reset, timer_0:reset_n]
	wire         rst_controller_003_reset_out_reset;                          // rst_controller_003:reset_out -> hps_emac_interface_splitter_0:rst_tx_n_o
	wire         hps_0_emac1_tx_reset_reset;                                  // hps_0:emac1_rst_clk_tx_n_o -> rst_controller_003:reset_in0
	wire         rst_controller_004_reset_out_reset;                          // rst_controller_004:reset_out -> mm_interconnect_0:hps_0_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset_reset
	wire         hps_0_h2f_reset_reset;                                       // hps_0:h2f_rst_n -> [rst_controller_004:reset_in0, rst_controller_005:reset_in0]
	wire         rst_controller_005_reset_out_reset;                          // rst_controller_005:reset_out -> mm_interconnect_1:hps_0_h2f_axi_master_agent_clk_reset_reset_bridge_in_reset_reset

	mn_soc_host_de10_nano_soc_hps_0 #(
		.F2S_Width (2),
		.S2F_Width (1)
	) hps_0 (
		.h2f_loan_in               (hps_0_h2f_loan_io_in),                                 //         h2f_loan_io.in
		.h2f_loan_out              (hps_0_h2f_loan_io_out),                                //                    .out
		.h2f_loan_oe               (hps_0_h2f_loan_io_oe),                                 //                    .oe
		.h2f_cold_rst_n            (hps_0_h2f_cold_reset_reset_n),                         //      h2f_cold_reset.reset_n
		.f2h_cold_rst_req_n        (hps_0_f2h_cold_reset_req_reset_n),                     //  f2h_cold_reset_req.reset_n
		.f2h_dbg_rst_req_n         (hps_0_f2h_debug_reset_req_reset_n),                    // f2h_debug_reset_req.reset_n
		.f2h_warm_rst_req_n        (hps_0_f2h_warm_reset_req_reset_n),                     //  f2h_warm_reset_req.reset_n
		.h2f_gp_in                 (hps_0_h2f_gp_gp_in),                                   //              h2f_gp.gp_in
		.h2f_gp_out                (hps_0_h2f_gp_gp_out),                                  //                    .gp_out
		.emac_ptp_ref_clk          (clk50_clk),                                            //  emac_ptp_ref_clock.clk
		.emac1_phy_txd_o           (hps_0_emac1_phy_txd_o),                                //               emac1.phy_txd_o
		.emac1_phy_txen_o          (hps_0_emac1_phy_txen_o),                               //                    .phy_txen_o
		.emac1_phy_txer_o          (hps_0_emac1_phy_txer_o),                               //                    .phy_txer_o
		.emac1_phy_rxdv_i          (hps_emac_interface_splitter_0_emac_phy_rxdv_i),        //                    .phy_rxdv_i
		.emac1_phy_rxer_i          (hps_emac_interface_splitter_0_emac_phy_rxer_i),        //                    .phy_rxer_i
		.emac1_phy_rxd_i           (hps_emac_interface_splitter_0_emac_phy_rxd_i),         //                    .phy_rxd_i
		.emac1_phy_col_i           (hps_emac_interface_splitter_0_emac_phy_col_i),         //                    .phy_col_i
		.emac1_phy_crs_i           (hps_emac_interface_splitter_0_emac_phy_crs_i),         //                    .phy_crs_i
		.emac1_gmii_mdo_o          (hps_0_emac1_gmii_mdo_o),                               //                    .gmii_mdo_o
		.emac1_gmii_mdo_o_e        (hps_0_emac1_gmii_mdo_o_e),                             //                    .gmii_mdo_o_e
		.emac1_gmii_mdi_i          (hps_emac_interface_splitter_0_emac_gmii_mdi_i),        //                    .gmii_mdi_i
		.emac1_ptp_pps_o           (hps_0_emac1_ptp_pps_o),                                //                    .ptp_pps_o
		.emac1_ptp_aux_ts_trig_i   (hps_emac_interface_splitter_0_emac_ptp_aux_ts_trig_i), //                    .ptp_aux_ts_trig_i
		.emac1_gmii_mdc_o          (hps_0_emac1_md_clk_clk),                               //        emac1_md_clk.clk
		.emac1_clk_rx_i            (hps_emac_interface_splitter_0_emac_rx_clk_in_clk),     //     emac1_rx_clk_in.clk
		.emac1_clk_tx_i            (hps_emac_interface_splitter_0_emac_tx_clk_in_clk),     //     emac1_tx_clk_in.clk
		.emac1_phy_txclk_o         (hps_0_emac1_gtx_clk_clk),                              //       emac1_gtx_clk.clk
		.emac1_rst_clk_tx_n_o      (hps_0_emac1_tx_reset_reset),                           //      emac1_tx_reset.reset_n
		.emac1_rst_clk_rx_n_o      (hps_0_emac1_rx_reset_reset),                           //      emac1_rx_reset.reset_n
		.mem_a                     (memory_mem_a),                                         //              memory.mem_a
		.mem_ba                    (memory_mem_ba),                                        //                    .mem_ba
		.mem_ck                    (memory_mem_ck),                                        //                    .mem_ck
		.mem_ck_n                  (memory_mem_ck_n),                                      //                    .mem_ck_n
		.mem_cke                   (memory_mem_cke),                                       //                    .mem_cke
		.mem_cs_n                  (memory_mem_cs_n),                                      //                    .mem_cs_n
		.mem_ras_n                 (memory_mem_ras_n),                                     //                    .mem_ras_n
		.mem_cas_n                 (memory_mem_cas_n),                                     //                    .mem_cas_n
		.mem_we_n                  (memory_mem_we_n),                                      //                    .mem_we_n
		.mem_reset_n               (memory_mem_reset_n),                                   //                    .mem_reset_n
		.mem_dq                    (memory_mem_dq),                                        //                    .mem_dq
		.mem_dqs                   (memory_mem_dqs),                                       //                    .mem_dqs
		.mem_dqs_n                 (memory_mem_dqs_n),                                     //                    .mem_dqs_n
		.mem_odt                   (memory_mem_odt),                                       //                    .mem_odt
		.mem_dm                    (memory_mem_dm),                                        //                    .mem_dm
		.oct_rzqin                 (memory_oct_rzqin),                                     //                    .oct_rzqin
		.hps_io_sdio_inst_CMD      (hps_0_hps_io_hps_io_sdio_inst_CMD),                    //              hps_io.hps_io_sdio_inst_CMD
		.hps_io_sdio_inst_D0       (hps_0_hps_io_hps_io_sdio_inst_D0),                     //                    .hps_io_sdio_inst_D0
		.hps_io_sdio_inst_D1       (hps_0_hps_io_hps_io_sdio_inst_D1),                     //                    .hps_io_sdio_inst_D1
		.hps_io_sdio_inst_CLK      (hps_0_hps_io_hps_io_sdio_inst_CLK),                    //                    .hps_io_sdio_inst_CLK
		.hps_io_sdio_inst_D2       (hps_0_hps_io_hps_io_sdio_inst_D2),                     //                    .hps_io_sdio_inst_D2
		.hps_io_sdio_inst_D3       (hps_0_hps_io_hps_io_sdio_inst_D3),                     //                    .hps_io_sdio_inst_D3
		.hps_io_usb1_inst_D0       (hps_0_hps_io_hps_io_usb1_inst_D0),                     //                    .hps_io_usb1_inst_D0
		.hps_io_usb1_inst_D1       (hps_0_hps_io_hps_io_usb1_inst_D1),                     //                    .hps_io_usb1_inst_D1
		.hps_io_usb1_inst_D2       (hps_0_hps_io_hps_io_usb1_inst_D2),                     //                    .hps_io_usb1_inst_D2
		.hps_io_usb1_inst_D3       (hps_0_hps_io_hps_io_usb1_inst_D3),                     //                    .hps_io_usb1_inst_D3
		.hps_io_usb1_inst_D4       (hps_0_hps_io_hps_io_usb1_inst_D4),                     //                    .hps_io_usb1_inst_D4
		.hps_io_usb1_inst_D5       (hps_0_hps_io_hps_io_usb1_inst_D5),                     //                    .hps_io_usb1_inst_D5
		.hps_io_usb1_inst_D6       (hps_0_hps_io_hps_io_usb1_inst_D6),                     //                    .hps_io_usb1_inst_D6
		.hps_io_usb1_inst_D7       (hps_0_hps_io_hps_io_usb1_inst_D7),                     //                    .hps_io_usb1_inst_D7
		.hps_io_usb1_inst_CLK      (hps_0_hps_io_hps_io_usb1_inst_CLK),                    //                    .hps_io_usb1_inst_CLK
		.hps_io_usb1_inst_STP      (hps_0_hps_io_hps_io_usb1_inst_STP),                    //                    .hps_io_usb1_inst_STP
		.hps_io_usb1_inst_DIR      (hps_0_hps_io_hps_io_usb1_inst_DIR),                    //                    .hps_io_usb1_inst_DIR
		.hps_io_usb1_inst_NXT      (hps_0_hps_io_hps_io_usb1_inst_NXT),                    //                    .hps_io_usb1_inst_NXT
		.hps_io_spim1_inst_CLK     (hps_0_hps_io_hps_io_spim1_inst_CLK),                   //                    .hps_io_spim1_inst_CLK
		.hps_io_spim1_inst_MOSI    (hps_0_hps_io_hps_io_spim1_inst_MOSI),                  //                    .hps_io_spim1_inst_MOSI
		.hps_io_spim1_inst_MISO    (hps_0_hps_io_hps_io_spim1_inst_MISO),                  //                    .hps_io_spim1_inst_MISO
		.hps_io_spim1_inst_SS0     (hps_0_hps_io_hps_io_spim1_inst_SS0),                   //                    .hps_io_spim1_inst_SS0
		.hps_io_uart0_inst_RX      (hps_0_hps_io_hps_io_uart0_inst_RX),                    //                    .hps_io_uart0_inst_RX
		.hps_io_uart0_inst_TX      (hps_0_hps_io_hps_io_uart0_inst_TX),                    //                    .hps_io_uart0_inst_TX
		.hps_io_i2c0_inst_SDA      (hps_0_hps_io_hps_io_i2c0_inst_SDA),                    //                    .hps_io_i2c0_inst_SDA
		.hps_io_i2c0_inst_SCL      (hps_0_hps_io_hps_io_i2c0_inst_SCL),                    //                    .hps_io_i2c0_inst_SCL
		.hps_io_i2c1_inst_SDA      (hps_0_hps_io_hps_io_i2c1_inst_SDA),                    //                    .hps_io_i2c1_inst_SDA
		.hps_io_i2c1_inst_SCL      (hps_0_hps_io_hps_io_i2c1_inst_SCL),                    //                    .hps_io_i2c1_inst_SCL
		.hps_io_gpio_inst_GPIO09   (hps_0_hps_io_hps_io_gpio_inst_GPIO09),                 //                    .hps_io_gpio_inst_GPIO09
		.hps_io_gpio_inst_GPIO35   (hps_0_hps_io_hps_io_gpio_inst_GPIO35),                 //                    .hps_io_gpio_inst_GPIO35
		.hps_io_gpio_inst_GPIO40   (hps_0_hps_io_hps_io_gpio_inst_GPIO40),                 //                    .hps_io_gpio_inst_GPIO40
		.hps_io_gpio_inst_GPIO53   (hps_0_hps_io_hps_io_gpio_inst_GPIO53),                 //                    .hps_io_gpio_inst_GPIO53
		.hps_io_gpio_inst_GPIO54   (hps_0_hps_io_hps_io_gpio_inst_GPIO54),                 //                    .hps_io_gpio_inst_GPIO54
		.hps_io_gpio_inst_GPIO61   (hps_0_hps_io_hps_io_gpio_inst_GPIO61),                 //                    .hps_io_gpio_inst_GPIO61
		.hps_io_gpio_inst_LOANIO20 (hps_0_hps_io_hps_io_gpio_inst_LOANIO20),               //                    .hps_io_gpio_inst_LOANIO20
		.hps_io_gpio_inst_LOANIO21 (hps_0_hps_io_hps_io_gpio_inst_LOANIO21),               //                    .hps_io_gpio_inst_LOANIO21
		.h2f_rst_n                 (hps_0_h2f_reset_reset),                                //           h2f_reset.reset_n
		.h2f_axi_clk               (clk100_clk),                                           //       h2f_axi_clock.clk
		.h2f_AWID                  (hps_0_h2f_axi_master_awid),                            //      h2f_axi_master.awid
		.h2f_AWADDR                (hps_0_h2f_axi_master_awaddr),                          //                    .awaddr
		.h2f_AWLEN                 (hps_0_h2f_axi_master_awlen),                           //                    .awlen
		.h2f_AWSIZE                (hps_0_h2f_axi_master_awsize),                          //                    .awsize
		.h2f_AWBURST               (hps_0_h2f_axi_master_awburst),                         //                    .awburst
		.h2f_AWLOCK                (hps_0_h2f_axi_master_awlock),                          //                    .awlock
		.h2f_AWCACHE               (hps_0_h2f_axi_master_awcache),                         //                    .awcache
		.h2f_AWPROT                (hps_0_h2f_axi_master_awprot),                          //                    .awprot
		.h2f_AWVALID               (hps_0_h2f_axi_master_awvalid),                         //                    .awvalid
		.h2f_AWREADY               (hps_0_h2f_axi_master_awready),                         //                    .awready
		.h2f_WID                   (hps_0_h2f_axi_master_wid),                             //                    .wid
		.h2f_WDATA                 (hps_0_h2f_axi_master_wdata),                           //                    .wdata
		.h2f_WSTRB                 (hps_0_h2f_axi_master_wstrb),                           //                    .wstrb
		.h2f_WLAST                 (hps_0_h2f_axi_master_wlast),                           //                    .wlast
		.h2f_WVALID                (hps_0_h2f_axi_master_wvalid),                          //                    .wvalid
		.h2f_WREADY                (hps_0_h2f_axi_master_wready),                          //                    .wready
		.h2f_BID                   (hps_0_h2f_axi_master_bid),                             //                    .bid
		.h2f_BRESP                 (hps_0_h2f_axi_master_bresp),                           //                    .bresp
		.h2f_BVALID                (hps_0_h2f_axi_master_bvalid),                          //                    .bvalid
		.h2f_BREADY                (hps_0_h2f_axi_master_bready),                          //                    .bready
		.h2f_ARID                  (hps_0_h2f_axi_master_arid),                            //                    .arid
		.h2f_ARADDR                (hps_0_h2f_axi_master_araddr),                          //                    .araddr
		.h2f_ARLEN                 (hps_0_h2f_axi_master_arlen),                           //                    .arlen
		.h2f_ARSIZE                (hps_0_h2f_axi_master_arsize),                          //                    .arsize
		.h2f_ARBURST               (hps_0_h2f_axi_master_arburst),                         //                    .arburst
		.h2f_ARLOCK                (hps_0_h2f_axi_master_arlock),                          //                    .arlock
		.h2f_ARCACHE               (hps_0_h2f_axi_master_arcache),                         //                    .arcache
		.h2f_ARPROT                (hps_0_h2f_axi_master_arprot),                          //                    .arprot
		.h2f_ARVALID               (hps_0_h2f_axi_master_arvalid),                         //                    .arvalid
		.h2f_ARREADY               (hps_0_h2f_axi_master_arready),                         //                    .arready
		.h2f_RID                   (hps_0_h2f_axi_master_rid),                             //                    .rid
		.h2f_RDATA                 (hps_0_h2f_axi_master_rdata),                           //                    .rdata
		.h2f_RRESP                 (hps_0_h2f_axi_master_rresp),                           //                    .rresp
		.h2f_RLAST                 (hps_0_h2f_axi_master_rlast),                           //                    .rlast
		.h2f_RVALID                (hps_0_h2f_axi_master_rvalid),                          //                    .rvalid
		.h2f_RREADY                (hps_0_h2f_axi_master_rready),                          //                    .rready
		.f2h_axi_clk               (clk50_clk),                                            //       f2h_axi_clock.clk
		.f2h_AWID                  (),                                                     //       f2h_axi_slave.awid
		.f2h_AWADDR                (),                                                     //                    .awaddr
		.f2h_AWLEN                 (),                                                     //                    .awlen
		.f2h_AWSIZE                (),                                                     //                    .awsize
		.f2h_AWBURST               (),                                                     //                    .awburst
		.f2h_AWLOCK                (),                                                     //                    .awlock
		.f2h_AWCACHE               (),                                                     //                    .awcache
		.f2h_AWPROT                (),                                                     //                    .awprot
		.f2h_AWVALID               (),                                                     //                    .awvalid
		.f2h_AWREADY               (),                                                     //                    .awready
		.f2h_AWUSER                (),                                                     //                    .awuser
		.f2h_WID                   (),                                                     //                    .wid
		.f2h_WDATA                 (),                                                     //                    .wdata
		.f2h_WSTRB                 (),                                                     //                    .wstrb
		.f2h_WLAST                 (),                                                     //                    .wlast
		.f2h_WVALID                (),                                                     //                    .wvalid
		.f2h_WREADY                (),                                                     //                    .wready
		.f2h_BID                   (),                                                     //                    .bid
		.f2h_BRESP                 (),                                                     //                    .bresp
		.f2h_BVALID                (),                                                     //                    .bvalid
		.f2h_BREADY                (),                                                     //                    .bready
		.f2h_ARID                  (),                                                     //                    .arid
		.f2h_ARADDR                (),                                                     //                    .araddr
		.f2h_ARLEN                 (),                                                     //                    .arlen
		.f2h_ARSIZE                (),                                                     //                    .arsize
		.f2h_ARBURST               (),                                                     //                    .arburst
		.f2h_ARLOCK                (),                                                     //                    .arlock
		.f2h_ARCACHE               (),                                                     //                    .arcache
		.f2h_ARPROT                (),                                                     //                    .arprot
		.f2h_ARVALID               (),                                                     //                    .arvalid
		.f2h_ARREADY               (),                                                     //                    .arready
		.f2h_ARUSER                (),                                                     //                    .aruser
		.f2h_RID                   (),                                                     //                    .rid
		.f2h_RDATA                 (),                                                     //                    .rdata
		.f2h_RRESP                 (),                                                     //                    .rresp
		.f2h_RLAST                 (),                                                     //                    .rlast
		.f2h_RVALID                (),                                                     //                    .rvalid
		.f2h_RREADY                (),                                                     //                    .rready
		.h2f_lw_axi_clk            (clk50_clk),                                            //    h2f_lw_axi_clock.clk
		.h2f_lw_AWID               (hps_0_h2f_lw_axi_master_awid),                         //   h2f_lw_axi_master.awid
		.h2f_lw_AWADDR             (hps_0_h2f_lw_axi_master_awaddr),                       //                    .awaddr
		.h2f_lw_AWLEN              (hps_0_h2f_lw_axi_master_awlen),                        //                    .awlen
		.h2f_lw_AWSIZE             (hps_0_h2f_lw_axi_master_awsize),                       //                    .awsize
		.h2f_lw_AWBURST            (hps_0_h2f_lw_axi_master_awburst),                      //                    .awburst
		.h2f_lw_AWLOCK             (hps_0_h2f_lw_axi_master_awlock),                       //                    .awlock
		.h2f_lw_AWCACHE            (hps_0_h2f_lw_axi_master_awcache),                      //                    .awcache
		.h2f_lw_AWPROT             (hps_0_h2f_lw_axi_master_awprot),                       //                    .awprot
		.h2f_lw_AWVALID            (hps_0_h2f_lw_axi_master_awvalid),                      //                    .awvalid
		.h2f_lw_AWREADY            (hps_0_h2f_lw_axi_master_awready),                      //                    .awready
		.h2f_lw_WID                (hps_0_h2f_lw_axi_master_wid),                          //                    .wid
		.h2f_lw_WDATA              (hps_0_h2f_lw_axi_master_wdata),                        //                    .wdata
		.h2f_lw_WSTRB              (hps_0_h2f_lw_axi_master_wstrb),                        //                    .wstrb
		.h2f_lw_WLAST              (hps_0_h2f_lw_axi_master_wlast),                        //                    .wlast
		.h2f_lw_WVALID             (hps_0_h2f_lw_axi_master_wvalid),                       //                    .wvalid
		.h2f_lw_WREADY             (hps_0_h2f_lw_axi_master_wready),                       //                    .wready
		.h2f_lw_BID                (hps_0_h2f_lw_axi_master_bid),                          //                    .bid
		.h2f_lw_BRESP              (hps_0_h2f_lw_axi_master_bresp),                        //                    .bresp
		.h2f_lw_BVALID             (hps_0_h2f_lw_axi_master_bvalid),                       //                    .bvalid
		.h2f_lw_BREADY             (hps_0_h2f_lw_axi_master_bready),                       //                    .bready
		.h2f_lw_ARID               (hps_0_h2f_lw_axi_master_arid),                         //                    .arid
		.h2f_lw_ARADDR             (hps_0_h2f_lw_axi_master_araddr),                       //                    .araddr
		.h2f_lw_ARLEN              (hps_0_h2f_lw_axi_master_arlen),                        //                    .arlen
		.h2f_lw_ARSIZE             (hps_0_h2f_lw_axi_master_arsize),                       //                    .arsize
		.h2f_lw_ARBURST            (hps_0_h2f_lw_axi_master_arburst),                      //                    .arburst
		.h2f_lw_ARLOCK             (hps_0_h2f_lw_axi_master_arlock),                       //                    .arlock
		.h2f_lw_ARCACHE            (hps_0_h2f_lw_axi_master_arcache),                      //                    .arcache
		.h2f_lw_ARPROT             (hps_0_h2f_lw_axi_master_arprot),                       //                    .arprot
		.h2f_lw_ARVALID            (hps_0_h2f_lw_axi_master_arvalid),                      //                    .arvalid
		.h2f_lw_ARREADY            (hps_0_h2f_lw_axi_master_arready),                      //                    .arready
		.h2f_lw_RID                (hps_0_h2f_lw_axi_master_rid),                          //                    .rid
		.h2f_lw_RDATA              (hps_0_h2f_lw_axi_master_rdata),                        //                    .rdata
		.h2f_lw_RRESP              (hps_0_h2f_lw_axi_master_rresp),                        //                    .rresp
		.h2f_lw_RLAST              (hps_0_h2f_lw_axi_master_rlast),                        //                    .rlast
		.h2f_lw_RVALID             (hps_0_h2f_lw_axi_master_rvalid),                       //                    .rvalid
		.h2f_lw_RREADY             (hps_0_h2f_lw_axi_master_rready),                       //                    .rready
		.f2h_irq_p0                (hps_0_f2h_irq0_irq),                                   //            f2h_irq0.irq
		.f2h_irq_p1                (hps_0_f2h_irq1_irq)                                    //            f2h_irq1.irq
	);

	mn_soc_host_de10_nano_soc_button_pio button_pio (
		.clk        (clk50_clk),                                  //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),            //               reset.reset_n
		.address    (mm_interconnect_0_button_pio_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_button_pio_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_button_pio_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_button_pio_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_button_pio_s1_readdata),   //                    .readdata
		.in_port    (button_pio_external_connection_export)       // external_connection.export
	);

	mn_soc_host_de10_nano_soc_dipsw_pio dipsw_pio (
		.clk        (clk50_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address    (mm_interconnect_0_dipsw_pio_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_dipsw_pio_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_dipsw_pio_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_dipsw_pio_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_dipsw_pio_s1_readdata),   //                    .readdata
		.in_port    (dipsw_pio_external_connection_export)       // external_connection.export
	);

	altera_avalon_mm_bridge #(
		.DATA_WIDTH        (32),
		.SYMBOL_WIDTH      (8),
		.HDL_ADDR_WIDTH    (27),
		.BURSTCOUNT_WIDTH  (1),
		.PIPELINE_COMMAND  (1),
		.PIPELINE_RESPONSE (1)
	) fpga_mem (
		.clk              (clk100_clk),                                  //   clk.clk
		.reset            (rst_controller_001_reset_out_reset),          // reset.reset
		.s0_waitrequest   (mm_interconnect_1_fpga_mem_s0_waitrequest),   //    s0.waitrequest
		.s0_readdata      (mm_interconnect_1_fpga_mem_s0_readdata),      //      .readdata
		.s0_readdatavalid (mm_interconnect_1_fpga_mem_s0_readdatavalid), //      .readdatavalid
		.s0_burstcount    (mm_interconnect_1_fpga_mem_s0_burstcount),    //      .burstcount
		.s0_writedata     (mm_interconnect_1_fpga_mem_s0_writedata),     //      .writedata
		.s0_address       (mm_interconnect_1_fpga_mem_s0_address),       //      .address
		.s0_write         (mm_interconnect_1_fpga_mem_s0_write),         //      .write
		.s0_read          (mm_interconnect_1_fpga_mem_s0_read),          //      .read
		.s0_byteenable    (mm_interconnect_1_fpga_mem_s0_byteenable),    //      .byteenable
		.s0_debugaccess   (mm_interconnect_1_fpga_mem_s0_debugaccess),   //      .debugaccess
		.m0_waitrequest   (fpga_mem_waitrequest),                        //    m0.waitrequest
		.m0_readdata      (fpga_mem_readdata),                           //      .readdata
		.m0_readdatavalid (fpga_mem_readdatavalid),                      //      .readdatavalid
		.m0_burstcount    (fpga_mem_burstcount),                         //      .burstcount
		.m0_writedata     (fpga_mem_writedata),                          //      .writedata
		.m0_address       (fpga_mem_address),                            //      .address
		.m0_write         (fpga_mem_write),                              //      .write
		.m0_read          (fpga_mem_read),                               //      .read
		.m0_byteenable    (fpga_mem_byteenable),                         //      .byteenable
		.m0_debugaccess   (fpga_mem_debugaccess)                         //      .debugaccess
	);

	altera_irq_bridge #(
		.IRQ_WIDTH (1)
	) hostif_irq (
		.clk          (clk50_clk),                          //          clk.clk
		.receiver_irq (hostif_irq_i_irq),                   // receiver_irq.irq
		.reset        (rst_controller_002_reset_out_reset), //    clk_reset.reset
		.sender0_irq  (irq_mapper_receiver0_irq),           //  sender0_irq.irq
		.sender1_irq  (),                                   //  (terminated)
		.sender2_irq  (),                                   //  (terminated)
		.sender3_irq  (),                                   //  (terminated)
		.sender4_irq  (),                                   //  (terminated)
		.sender5_irq  (),                                   //  (terminated)
		.sender6_irq  (),                                   //  (terminated)
		.sender7_irq  (),                                   //  (terminated)
		.sender8_irq  (),                                   //  (terminated)
		.sender9_irq  (),                                   //  (terminated)
		.sender10_irq (),                                   //  (terminated)
		.sender11_irq (),                                   //  (terminated)
		.sender12_irq (),                                   //  (terminated)
		.sender13_irq (),                                   //  (terminated)
		.sender14_irq (),                                   //  (terminated)
		.sender15_irq (),                                   //  (terminated)
		.sender16_irq (),                                   //  (terminated)
		.sender17_irq (),                                   //  (terminated)
		.sender18_irq (),                                   //  (terminated)
		.sender19_irq (),                                   //  (terminated)
		.sender20_irq (),                                   //  (terminated)
		.sender21_irq (),                                   //  (terminated)
		.sender22_irq (),                                   //  (terminated)
		.sender23_irq (),                                   //  (terminated)
		.sender24_irq (),                                   //  (terminated)
		.sender25_irq (),                                   //  (terminated)
		.sender26_irq (),                                   //  (terminated)
		.sender27_irq (),                                   //  (terminated)
		.sender28_irq (),                                   //  (terminated)
		.sender29_irq (),                                   //  (terminated)
		.sender30_irq (),                                   //  (terminated)
		.sender31_irq ()                                    //  (terminated)
	);

	altera_avalon_mm_bridge #(
		.DATA_WIDTH        (32),
		.SYMBOL_WIDTH      (8),
		.HDL_ADDR_WIDTH    (18),
		.BURSTCOUNT_WIDTH  (1),
		.PIPELINE_COMMAND  (1),
		.PIPELINE_RESPONSE (1)
	) lw_bridge (
		.clk              (clk50_clk),                                    //   clk.clk
		.reset            (rst_controller_002_reset_out_reset),           // reset.reset
		.s0_waitrequest   (mm_interconnect_0_lw_bridge_s0_waitrequest),   //    s0.waitrequest
		.s0_readdata      (mm_interconnect_0_lw_bridge_s0_readdata),      //      .readdata
		.s0_readdatavalid (mm_interconnect_0_lw_bridge_s0_readdatavalid), //      .readdatavalid
		.s0_burstcount    (mm_interconnect_0_lw_bridge_s0_burstcount),    //      .burstcount
		.s0_writedata     (mm_interconnect_0_lw_bridge_s0_writedata),     //      .writedata
		.s0_address       (mm_interconnect_0_lw_bridge_s0_address),       //      .address
		.s0_write         (mm_interconnect_0_lw_bridge_s0_write),         //      .write
		.s0_read          (mm_interconnect_0_lw_bridge_s0_read),          //      .read
		.s0_byteenable    (mm_interconnect_0_lw_bridge_s0_byteenable),    //      .byteenable
		.s0_debugaccess   (mm_interconnect_0_lw_bridge_s0_debugaccess),   //      .debugaccess
		.m0_waitrequest   (lw_bridge_m0_waitrequest),                     //    m0.waitrequest
		.m0_readdata      (lw_bridge_m0_readdata),                        //      .readdata
		.m0_readdatavalid (lw_bridge_m0_readdatavalid),                   //      .readdatavalid
		.m0_burstcount    (lw_bridge_m0_burstcount),                      //      .burstcount
		.m0_writedata     (lw_bridge_m0_writedata),                       //      .writedata
		.m0_address       (lw_bridge_m0_address),                         //      .address
		.m0_write         (lw_bridge_m0_write),                           //      .write
		.m0_read          (lw_bridge_m0_read),                            //      .read
		.m0_byteenable    (lw_bridge_m0_byteenable),                      //      .byteenable
		.m0_debugaccess   (lw_bridge_m0_debugaccess)                      //      .debugaccess
	);

	mn_soc_host_de10_nano_soc_jtag_uart_0 jtag_uart_0 (
		.clk            (clk50_clk),                                                   //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                             //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver1_irq)                                     //               irq.irq
	);

	mn_soc_host_de10_nano_soc_timer_0 timer_0 (
		.clk        (clk50_clk),                               //   clk.clk
		.reset_n    (~rst_controller_002_reset_out_reset),     // reset.reset_n
		.address    (mm_interconnect_0_timer_0_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer_0_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer_0_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer_0_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer_0_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver2_irq)                 //   irq.irq
	);

	altera_hps_emac_interface_splitter #(
		.MAC_SPEED_CSR_ENABLE (1)
	) hps_emac_interface_splitter_0 (
		.phy_txclk_o        (hps_0_emac1_gtx_clk_clk),                                //   emac_gtx_clk.clk
		.clk_tx_i           (hps_emac_interface_splitter_0_emac_tx_clk_in_clk),       // emac_tx_clk_in.clk
		.clk_rx_i           (hps_emac_interface_splitter_0_emac_rx_clk_in_clk),       // emac_rx_clk_in.clk
		.rst_tx_n_o         (~rst_controller_003_reset_out_reset),                    //  emac_tx_reset.reset_n
		.rst_rx_n_o         (hps_0_emac1_rx_reset_reset),                             //  emac_rx_reset.reset_n
		.mac_tx_clk_i       (hps_emac_interface_splitter_0_hps_gmii_phy_tx_clk_i),    //       hps_gmii.phy_tx_clk_i
		.mac_rx_clk         (hps_emac_interface_splitter_0_hps_gmii_phy_rx_clk_i),    //               .phy_rx_clk_i
		.mac_rxdv           (hps_emac_interface_splitter_0_hps_gmii_phy_rxdv_i),      //               .phy_rxdv_i
		.mac_rxer           (hps_emac_interface_splitter_0_hps_gmii_phy_rxer_i),      //               .phy_rxer_i
		.mac_rxd            (hps_emac_interface_splitter_0_hps_gmii_phy_rxd_i),       //               .phy_rxd_i
		.mac_col            (hps_emac_interface_splitter_0_hps_gmii_phy_col_i),       //               .phy_col_i
		.mac_crs            (hps_emac_interface_splitter_0_hps_gmii_phy_crs_i),       //               .phy_crs_i
		.mac_tx_clk_o       (hps_emac_interface_splitter_0_hps_gmii_phy_tx_clk_o),    //               .phy_tx_clk_o
		.mac_rst_tx_n       (hps_emac_interface_splitter_0_hps_gmii_rst_tx_n),        //               .rst_tx_n
		.mac_rst_rx_n       (hps_emac_interface_splitter_0_hps_gmii_rst_rx_n),        //               .rst_rx_n
		.mac_txd            (hps_emac_interface_splitter_0_hps_gmii_phy_txd_o),       //               .phy_txd_o
		.mac_txen           (hps_emac_interface_splitter_0_hps_gmii_phy_txen_o),      //               .phy_txen_o
		.mac_txer           (hps_emac_interface_splitter_0_hps_gmii_phy_txer_o),      //               .phy_txer_o
		.mac_speed          (hps_emac_interface_splitter_0_hps_gmii_phy_mac_speed_o), //               .phy_mac_speed_o
		.mdi_in             (hps_emac_interface_splitter_0_mdio_gmii_mdi_i),          //           mdio.gmii_mdi_i
		.mdo_out            (hps_emac_interface_splitter_0_mdio_gmii_mdo_o),          //               .gmii_mdo_o
		.mdo_out_en         (hps_emac_interface_splitter_0_mdio_gmii_mdo_o_e),        //               .gmii_mdo_o_e
		.ptp_aux_ts_trig_in (hps_emac_interface_splitter_0_ptp_ptp_aux_ts_trig_i),    //            ptp.ptp_aux_ts_trig_i
		.ptp_pps_out        (hps_emac_interface_splitter_0_ptp_ptp_pps_o),            //               .ptp_pps_o
		.clk                (clk50_clk),                                              //     peri_clock.clk
		.rst_n              (~rst_controller_reset_out_reset),                        //     peri_reset.reset_n
		.read               (),                                                       //   avalon_slave.read
		.write              (),                                                       //               .write
		.writedata          (),                                                       //               .writedata
		.readdata           (),                                                       //               .readdata
		.addr               (),                                                       //               .address
		.phy_txd_o          (hps_0_emac1_phy_txd_o),                                  //           emac.phy_txd_o
		.phy_txen_o         (hps_0_emac1_phy_txen_o),                                 //               .phy_txen_o
		.phy_txer_o         (hps_0_emac1_phy_txer_o),                                 //               .phy_txer_o
		.mdo_o              (hps_0_emac1_gmii_mdo_o),                                 //               .gmii_mdo_o
		.mdo_o_e            (hps_0_emac1_gmii_mdo_o_e),                               //               .gmii_mdo_o_e
		.ptp_pps_o          (hps_0_emac1_ptp_pps_o),                                  //               .ptp_pps_o
		.phy_rxdv_i         (hps_emac_interface_splitter_0_emac_phy_rxdv_i),          //               .phy_rxdv_i
		.phy_rxer_i         (hps_emac_interface_splitter_0_emac_phy_rxer_i),          //               .phy_rxer_i
		.phy_rxd_i          (hps_emac_interface_splitter_0_emac_phy_rxd_i),           //               .phy_rxd_i
		.phy_col_i          (hps_emac_interface_splitter_0_emac_phy_col_i),           //               .phy_col_i
		.phy_crs_i          (hps_emac_interface_splitter_0_emac_phy_crs_i),           //               .phy_crs_i
		.mdi_i              (hps_emac_interface_splitter_0_emac_gmii_mdi_i),          //               .gmii_mdi_i
		.ptp_aux_ts_trig_i  (hps_emac_interface_splitter_0_emac_ptp_aux_ts_trig_i),   //               .ptp_aux_ts_trig_i
		.phy_mac_speed_o    (2'b00)                                                   //    (terminated)
	);

	mn_soc_host_de10_nano_soc_mm_interconnect_0 mm_interconnect_0 (
		.hps_0_h2f_lw_axi_master_awid                                        (hps_0_h2f_lw_axi_master_awid),                                //                                       hps_0_h2f_lw_axi_master.awid
		.hps_0_h2f_lw_axi_master_awaddr                                      (hps_0_h2f_lw_axi_master_awaddr),                              //                                                              .awaddr
		.hps_0_h2f_lw_axi_master_awlen                                       (hps_0_h2f_lw_axi_master_awlen),                               //                                                              .awlen
		.hps_0_h2f_lw_axi_master_awsize                                      (hps_0_h2f_lw_axi_master_awsize),                              //                                                              .awsize
		.hps_0_h2f_lw_axi_master_awburst                                     (hps_0_h2f_lw_axi_master_awburst),                             //                                                              .awburst
		.hps_0_h2f_lw_axi_master_awlock                                      (hps_0_h2f_lw_axi_master_awlock),                              //                                                              .awlock
		.hps_0_h2f_lw_axi_master_awcache                                     (hps_0_h2f_lw_axi_master_awcache),                             //                                                              .awcache
		.hps_0_h2f_lw_axi_master_awprot                                      (hps_0_h2f_lw_axi_master_awprot),                              //                                                              .awprot
		.hps_0_h2f_lw_axi_master_awvalid                                     (hps_0_h2f_lw_axi_master_awvalid),                             //                                                              .awvalid
		.hps_0_h2f_lw_axi_master_awready                                     (hps_0_h2f_lw_axi_master_awready),                             //                                                              .awready
		.hps_0_h2f_lw_axi_master_wid                                         (hps_0_h2f_lw_axi_master_wid),                                 //                                                              .wid
		.hps_0_h2f_lw_axi_master_wdata                                       (hps_0_h2f_lw_axi_master_wdata),                               //                                                              .wdata
		.hps_0_h2f_lw_axi_master_wstrb                                       (hps_0_h2f_lw_axi_master_wstrb),                               //                                                              .wstrb
		.hps_0_h2f_lw_axi_master_wlast                                       (hps_0_h2f_lw_axi_master_wlast),                               //                                                              .wlast
		.hps_0_h2f_lw_axi_master_wvalid                                      (hps_0_h2f_lw_axi_master_wvalid),                              //                                                              .wvalid
		.hps_0_h2f_lw_axi_master_wready                                      (hps_0_h2f_lw_axi_master_wready),                              //                                                              .wready
		.hps_0_h2f_lw_axi_master_bid                                         (hps_0_h2f_lw_axi_master_bid),                                 //                                                              .bid
		.hps_0_h2f_lw_axi_master_bresp                                       (hps_0_h2f_lw_axi_master_bresp),                               //                                                              .bresp
		.hps_0_h2f_lw_axi_master_bvalid                                      (hps_0_h2f_lw_axi_master_bvalid),                              //                                                              .bvalid
		.hps_0_h2f_lw_axi_master_bready                                      (hps_0_h2f_lw_axi_master_bready),                              //                                                              .bready
		.hps_0_h2f_lw_axi_master_arid                                        (hps_0_h2f_lw_axi_master_arid),                                //                                                              .arid
		.hps_0_h2f_lw_axi_master_araddr                                      (hps_0_h2f_lw_axi_master_araddr),                              //                                                              .araddr
		.hps_0_h2f_lw_axi_master_arlen                                       (hps_0_h2f_lw_axi_master_arlen),                               //                                                              .arlen
		.hps_0_h2f_lw_axi_master_arsize                                      (hps_0_h2f_lw_axi_master_arsize),                              //                                                              .arsize
		.hps_0_h2f_lw_axi_master_arburst                                     (hps_0_h2f_lw_axi_master_arburst),                             //                                                              .arburst
		.hps_0_h2f_lw_axi_master_arlock                                      (hps_0_h2f_lw_axi_master_arlock),                              //                                                              .arlock
		.hps_0_h2f_lw_axi_master_arcache                                     (hps_0_h2f_lw_axi_master_arcache),                             //                                                              .arcache
		.hps_0_h2f_lw_axi_master_arprot                                      (hps_0_h2f_lw_axi_master_arprot),                              //                                                              .arprot
		.hps_0_h2f_lw_axi_master_arvalid                                     (hps_0_h2f_lw_axi_master_arvalid),                             //                                                              .arvalid
		.hps_0_h2f_lw_axi_master_arready                                     (hps_0_h2f_lw_axi_master_arready),                             //                                                              .arready
		.hps_0_h2f_lw_axi_master_rid                                         (hps_0_h2f_lw_axi_master_rid),                                 //                                                              .rid
		.hps_0_h2f_lw_axi_master_rdata                                       (hps_0_h2f_lw_axi_master_rdata),                               //                                                              .rdata
		.hps_0_h2f_lw_axi_master_rresp                                       (hps_0_h2f_lw_axi_master_rresp),                               //                                                              .rresp
		.hps_0_h2f_lw_axi_master_rlast                                       (hps_0_h2f_lw_axi_master_rlast),                               //                                                              .rlast
		.hps_0_h2f_lw_axi_master_rvalid                                      (hps_0_h2f_lw_axi_master_rvalid),                              //                                                              .rvalid
		.hps_0_h2f_lw_axi_master_rready                                      (hps_0_h2f_lw_axi_master_rready),                              //                                                              .rready
		.clk_50_clk_clk                                                      (clk50_clk),                                                   //                                                    clk_50_clk.clk
		.dipsw_pio_reset_reset_bridge_in_reset_reset                         (rst_controller_reset_out_reset),                              //                         dipsw_pio_reset_reset_bridge_in_reset.reset
		.hps_0_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset_reset (rst_controller_004_reset_out_reset),                          // hps_0_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset.reset
		.lw_bridge_reset_reset_bridge_in_reset_reset                         (rst_controller_002_reset_out_reset),                          //                         lw_bridge_reset_reset_bridge_in_reset.reset
		.button_pio_s1_address                                               (mm_interconnect_0_button_pio_s1_address),                     //                                                 button_pio_s1.address
		.button_pio_s1_write                                                 (mm_interconnect_0_button_pio_s1_write),                       //                                                              .write
		.button_pio_s1_readdata                                              (mm_interconnect_0_button_pio_s1_readdata),                    //                                                              .readdata
		.button_pio_s1_writedata                                             (mm_interconnect_0_button_pio_s1_writedata),                   //                                                              .writedata
		.button_pio_s1_chipselect                                            (mm_interconnect_0_button_pio_s1_chipselect),                  //                                                              .chipselect
		.dipsw_pio_s1_address                                                (mm_interconnect_0_dipsw_pio_s1_address),                      //                                                  dipsw_pio_s1.address
		.dipsw_pio_s1_write                                                  (mm_interconnect_0_dipsw_pio_s1_write),                        //                                                              .write
		.dipsw_pio_s1_readdata                                               (mm_interconnect_0_dipsw_pio_s1_readdata),                     //                                                              .readdata
		.dipsw_pio_s1_writedata                                              (mm_interconnect_0_dipsw_pio_s1_writedata),                    //                                                              .writedata
		.dipsw_pio_s1_chipselect                                             (mm_interconnect_0_dipsw_pio_s1_chipselect),                   //                                                              .chipselect
		.jtag_uart_0_avalon_jtag_slave_address                               (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),     //                                 jtag_uart_0_avalon_jtag_slave.address
		.jtag_uart_0_avalon_jtag_slave_write                                 (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),       //                                                              .write
		.jtag_uart_0_avalon_jtag_slave_read                                  (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),        //                                                              .read
		.jtag_uart_0_avalon_jtag_slave_readdata                              (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),    //                                                              .readdata
		.jtag_uart_0_avalon_jtag_slave_writedata                             (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),   //                                                              .writedata
		.jtag_uart_0_avalon_jtag_slave_waitrequest                           (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest), //                                                              .waitrequest
		.jtag_uart_0_avalon_jtag_slave_chipselect                            (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),  //                                                              .chipselect
		.lw_bridge_s0_address                                                (mm_interconnect_0_lw_bridge_s0_address),                      //                                                  lw_bridge_s0.address
		.lw_bridge_s0_write                                                  (mm_interconnect_0_lw_bridge_s0_write),                        //                                                              .write
		.lw_bridge_s0_read                                                   (mm_interconnect_0_lw_bridge_s0_read),                         //                                                              .read
		.lw_bridge_s0_readdata                                               (mm_interconnect_0_lw_bridge_s0_readdata),                     //                                                              .readdata
		.lw_bridge_s0_writedata                                              (mm_interconnect_0_lw_bridge_s0_writedata),                    //                                                              .writedata
		.lw_bridge_s0_burstcount                                             (mm_interconnect_0_lw_bridge_s0_burstcount),                   //                                                              .burstcount
		.lw_bridge_s0_byteenable                                             (mm_interconnect_0_lw_bridge_s0_byteenable),                   //                                                              .byteenable
		.lw_bridge_s0_readdatavalid                                          (mm_interconnect_0_lw_bridge_s0_readdatavalid),                //                                                              .readdatavalid
		.lw_bridge_s0_waitrequest                                            (mm_interconnect_0_lw_bridge_s0_waitrequest),                  //                                                              .waitrequest
		.lw_bridge_s0_debugaccess                                            (mm_interconnect_0_lw_bridge_s0_debugaccess),                  //                                                              .debugaccess
		.timer_0_s1_address                                                  (mm_interconnect_0_timer_0_s1_address),                        //                                                    timer_0_s1.address
		.timer_0_s1_write                                                    (mm_interconnect_0_timer_0_s1_write),                          //                                                              .write
		.timer_0_s1_readdata                                                 (mm_interconnect_0_timer_0_s1_readdata),                       //                                                              .readdata
		.timer_0_s1_writedata                                                (mm_interconnect_0_timer_0_s1_writedata),                      //                                                              .writedata
		.timer_0_s1_chipselect                                               (mm_interconnect_0_timer_0_s1_chipselect)                      //                                                              .chipselect
	);

	mn_soc_host_de10_nano_soc_mm_interconnect_1 mm_interconnect_1 (
		.hps_0_h2f_axi_master_awid                                        (hps_0_h2f_axi_master_awid),                   //                                       hps_0_h2f_axi_master.awid
		.hps_0_h2f_axi_master_awaddr                                      (hps_0_h2f_axi_master_awaddr),                 //                                                           .awaddr
		.hps_0_h2f_axi_master_awlen                                       (hps_0_h2f_axi_master_awlen),                  //                                                           .awlen
		.hps_0_h2f_axi_master_awsize                                      (hps_0_h2f_axi_master_awsize),                 //                                                           .awsize
		.hps_0_h2f_axi_master_awburst                                     (hps_0_h2f_axi_master_awburst),                //                                                           .awburst
		.hps_0_h2f_axi_master_awlock                                      (hps_0_h2f_axi_master_awlock),                 //                                                           .awlock
		.hps_0_h2f_axi_master_awcache                                     (hps_0_h2f_axi_master_awcache),                //                                                           .awcache
		.hps_0_h2f_axi_master_awprot                                      (hps_0_h2f_axi_master_awprot),                 //                                                           .awprot
		.hps_0_h2f_axi_master_awvalid                                     (hps_0_h2f_axi_master_awvalid),                //                                                           .awvalid
		.hps_0_h2f_axi_master_awready                                     (hps_0_h2f_axi_master_awready),                //                                                           .awready
		.hps_0_h2f_axi_master_wid                                         (hps_0_h2f_axi_master_wid),                    //                                                           .wid
		.hps_0_h2f_axi_master_wdata                                       (hps_0_h2f_axi_master_wdata),                  //                                                           .wdata
		.hps_0_h2f_axi_master_wstrb                                       (hps_0_h2f_axi_master_wstrb),                  //                                                           .wstrb
		.hps_0_h2f_axi_master_wlast                                       (hps_0_h2f_axi_master_wlast),                  //                                                           .wlast
		.hps_0_h2f_axi_master_wvalid                                      (hps_0_h2f_axi_master_wvalid),                 //                                                           .wvalid
		.hps_0_h2f_axi_master_wready                                      (hps_0_h2f_axi_master_wready),                 //                                                           .wready
		.hps_0_h2f_axi_master_bid                                         (hps_0_h2f_axi_master_bid),                    //                                                           .bid
		.hps_0_h2f_axi_master_bresp                                       (hps_0_h2f_axi_master_bresp),                  //                                                           .bresp
		.hps_0_h2f_axi_master_bvalid                                      (hps_0_h2f_axi_master_bvalid),                 //                                                           .bvalid
		.hps_0_h2f_axi_master_bready                                      (hps_0_h2f_axi_master_bready),                 //                                                           .bready
		.hps_0_h2f_axi_master_arid                                        (hps_0_h2f_axi_master_arid),                   //                                                           .arid
		.hps_0_h2f_axi_master_araddr                                      (hps_0_h2f_axi_master_araddr),                 //                                                           .araddr
		.hps_0_h2f_axi_master_arlen                                       (hps_0_h2f_axi_master_arlen),                  //                                                           .arlen
		.hps_0_h2f_axi_master_arsize                                      (hps_0_h2f_axi_master_arsize),                 //                                                           .arsize
		.hps_0_h2f_axi_master_arburst                                     (hps_0_h2f_axi_master_arburst),                //                                                           .arburst
		.hps_0_h2f_axi_master_arlock                                      (hps_0_h2f_axi_master_arlock),                 //                                                           .arlock
		.hps_0_h2f_axi_master_arcache                                     (hps_0_h2f_axi_master_arcache),                //                                                           .arcache
		.hps_0_h2f_axi_master_arprot                                      (hps_0_h2f_axi_master_arprot),                 //                                                           .arprot
		.hps_0_h2f_axi_master_arvalid                                     (hps_0_h2f_axi_master_arvalid),                //                                                           .arvalid
		.hps_0_h2f_axi_master_arready                                     (hps_0_h2f_axi_master_arready),                //                                                           .arready
		.hps_0_h2f_axi_master_rid                                         (hps_0_h2f_axi_master_rid),                    //                                                           .rid
		.hps_0_h2f_axi_master_rdata                                       (hps_0_h2f_axi_master_rdata),                  //                                                           .rdata
		.hps_0_h2f_axi_master_rresp                                       (hps_0_h2f_axi_master_rresp),                  //                                                           .rresp
		.hps_0_h2f_axi_master_rlast                                       (hps_0_h2f_axi_master_rlast),                  //                                                           .rlast
		.hps_0_h2f_axi_master_rvalid                                      (hps_0_h2f_axi_master_rvalid),                 //                                                           .rvalid
		.hps_0_h2f_axi_master_rready                                      (hps_0_h2f_axi_master_rready),                 //                                                           .rready
		.clk_100_clk_clk                                                  (clk100_clk),                                  //                                                clk_100_clk.clk
		.fpga_mem_reset_reset_bridge_in_reset_reset                       (rst_controller_001_reset_out_reset),          //                       fpga_mem_reset_reset_bridge_in_reset.reset
		.hps_0_h2f_axi_master_agent_clk_reset_reset_bridge_in_reset_reset (rst_controller_005_reset_out_reset),          // hps_0_h2f_axi_master_agent_clk_reset_reset_bridge_in_reset.reset
		.fpga_mem_s0_address                                              (mm_interconnect_1_fpga_mem_s0_address),       //                                                fpga_mem_s0.address
		.fpga_mem_s0_write                                                (mm_interconnect_1_fpga_mem_s0_write),         //                                                           .write
		.fpga_mem_s0_read                                                 (mm_interconnect_1_fpga_mem_s0_read),          //                                                           .read
		.fpga_mem_s0_readdata                                             (mm_interconnect_1_fpga_mem_s0_readdata),      //                                                           .readdata
		.fpga_mem_s0_writedata                                            (mm_interconnect_1_fpga_mem_s0_writedata),     //                                                           .writedata
		.fpga_mem_s0_burstcount                                           (mm_interconnect_1_fpga_mem_s0_burstcount),    //                                                           .burstcount
		.fpga_mem_s0_byteenable                                           (mm_interconnect_1_fpga_mem_s0_byteenable),    //                                                           .byteenable
		.fpga_mem_s0_readdatavalid                                        (mm_interconnect_1_fpga_mem_s0_readdatavalid), //                                                           .readdatavalid
		.fpga_mem_s0_waitrequest                                          (mm_interconnect_1_fpga_mem_s0_waitrequest),   //                                                           .waitrequest
		.fpga_mem_s0_debugaccess                                          (mm_interconnect_1_fpga_mem_s0_debugaccess)    //                                                           .debugaccess
	);

	mn_soc_host_de10_nano_soc_irq_mapper irq_mapper (
		.clk           (),                         //       clk.clk
		.reset         (),                         // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq), // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq), // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq), // receiver2.irq
		.sender_irq    (hps_0_f2h_irq0_irq)        //    sender.irq
	);

	mn_soc_host_de10_nano_soc_irq_mapper_001 irq_mapper_001 (
		.clk        (),                   //       clk.clk
		.reset      (),                   // clk_reset.reset
		.sender_irq (hps_0_f2h_irq1_irq)  //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_clk50_reset_n),           // reset_in0.reset
		.clk            (clk50_clk),                      //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_clk50_reset_n),               // reset_in0.reset
		.clk            (clk100_clk),                         //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_002 (
		.reset_in0      (~reset_clk100_reset_n),              // reset_in0.reset
		.reset_in1      (~reset_clk50_reset_n),               // reset_in1.reset
		.clk            (clk50_clk),                          //       clk.clk
		.reset_out      (rst_controller_002_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_003 (
		.reset_in0      (~hps_0_emac1_tx_reset_reset),        // reset_in0.reset
		.clk            (hps_0_emac1_gtx_clk_clk),            //       clk.clk
		.reset_out      (rst_controller_003_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_004 (
		.reset_in0      (~hps_0_h2f_reset_reset),             // reset_in0.reset
		.clk            (clk50_clk),                          //       clk.clk
		.reset_out      (rst_controller_004_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_005 (
		.reset_in0      (~hps_0_h2f_reset_reset),             // reset_in0.reset
		.clk            (clk100_clk),                         //       clk.clk
		.reset_out      (rst_controller_005_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
