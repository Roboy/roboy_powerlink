// soc_system_pcp_0.v

// Generated using ACDS version 14.0 200 at 2018.02.08.18:46:03

`timescale 1 ps / 1 ps
module soc_system_pcp_0 (
		input  wire        clk50_clk,                                //                             clk50.clk
		input  wire        rst_clk50_reset_n,                        //                         rst_clk50.reset_n
		input  wire        clk100_clk,                               //                            clk100.clk
		input  wire        rst_clk100_reset_n,                       //                        rst_clk100.reset_n
		output wire [7:0]  benchmark_pio_external_connection_export, // benchmark_pio_external_connection.export
		input  wire        slow_bridge_waitrequest,                  //                       slow_bridge.waitrequest
		input  wire [31:0] slow_bridge_readdata,                     //                                  .readdata
		input  wire        slow_bridge_readdatavalid,                //                                  .readdatavalid
		output wire [0:0]  slow_bridge_burstcount,                   //                                  .burstcount
		output wire [31:0] slow_bridge_writedata,                    //                                  .writedata
		output wire [18:0] slow_bridge_address,                      //                                  .address
		output wire        slow_bridge_write,                        //                                  .write
		output wire        slow_bridge_read,                         //                                  .read
		output wire [3:0]  slow_bridge_byteenable,                   //                                  .byteenable
		output wire        slow_bridge_debugaccess,                  //                                  .debugaccess
		input  wire        cpu_bridge_waitrequest,                   //                        cpu_bridge.waitrequest
		input  wire [31:0] cpu_bridge_readdata,                      //                                  .readdata
		input  wire        cpu_bridge_readdatavalid,                 //                                  .readdatavalid
		output wire [0:0]  cpu_bridge_burstcount,                    //                                  .burstcount
		output wire [31:0] cpu_bridge_writedata,                     //                                  .writedata
		output wire [21:0] cpu_bridge_address,                       //                                  .address
		output wire        cpu_bridge_write,                         //                                  .write
		output wire        cpu_bridge_read,                          //                                  .read
		output wire [3:0]  cpu_bridge_byteenable,                    //                                  .byteenable
		output wire        cpu_bridge_debugaccess,                   //                                  .debugaccess
		input  wire [0:0]  sync_irq_irq,                             //                          sync_irq.irq
		input  wire [0:0]  mac_irq_irq,                              //                           mac_irq.irq
		input  wire        flash_bridge_waitrequest,                 //                      flash_bridge.waitrequest
		input  wire [31:0] flash_bridge_readdata,                    //                                  .readdata
		input  wire        flash_bridge_readdatavalid,               //                                  .readdatavalid
		output wire [0:0]  flash_bridge_burstcount,                  //                                  .burstcount
		output wire [31:0] flash_bridge_writedata,                   //                                  .writedata
		output wire [21:0] flash_bridge_address,                     //                                  .address
		output wire        flash_bridge_write,                       //                                  .write
		output wire        flash_bridge_read,                        //                                  .read
		output wire [3:0]  flash_bridge_byteenable,                  //                                  .byteenable
		output wire        flash_bridge_debugaccess,                 //                                  .debugaccess
		input  wire [3:0]  gp_irq_irq,                               //                            gp_irq.irq
		input  wire        cpu_resetrequest_resetrequest,            //                  cpu_resetrequest.resetrequest
		output wire        cpu_resetrequest_resettaken,              //                                  .resettaken
		output wire        jtag_reset_reset,                         //                        jtag_reset.reset
		output wire [1:0]  powerlink_led_export                      //                     powerlink_led.export
	);

	wire         cpu_0_instruction_master_waitrequest;                        // mm_interconnect_0:cpu_0_instruction_master_waitrequest -> cpu_0:i_waitrequest
	wire  [25:0] cpu_0_instruction_master_address;                            // cpu_0:i_address -> mm_interconnect_0:cpu_0_instruction_master_address
	wire         cpu_0_instruction_master_read;                               // cpu_0:i_read -> mm_interconnect_0:cpu_0_instruction_master_read
	wire  [31:0] cpu_0_instruction_master_readdata;                           // mm_interconnect_0:cpu_0_instruction_master_readdata -> cpu_0:i_readdata
	wire         cpu_0_instruction_master_readdatavalid;                      // mm_interconnect_0:cpu_0_instruction_master_readdatavalid -> cpu_0:i_readdatavalid
	wire         cpu_0_data_master_waitrequest;                               // mm_interconnect_0:cpu_0_data_master_waitrequest -> cpu_0:d_waitrequest
	wire  [31:0] cpu_0_data_master_writedata;                                 // cpu_0:d_writedata -> mm_interconnect_0:cpu_0_data_master_writedata
	wire  [29:0] cpu_0_data_master_address;                                   // cpu_0:d_address -> mm_interconnect_0:cpu_0_data_master_address
	wire         cpu_0_data_master_write;                                     // cpu_0:d_write -> mm_interconnect_0:cpu_0_data_master_write
	wire         cpu_0_data_master_read;                                      // cpu_0:d_read -> mm_interconnect_0:cpu_0_data_master_read
	wire  [31:0] cpu_0_data_master_readdata;                                  // mm_interconnect_0:cpu_0_data_master_readdata -> cpu_0:d_readdata
	wire         cpu_0_data_master_debugaccess;                               // cpu_0:jtag_debug_module_debugaccess_to_roms -> mm_interconnect_0:cpu_0_data_master_debugaccess
	wire   [3:0] cpu_0_data_master_byteenable;                                // cpu_0:d_byteenable -> mm_interconnect_0:cpu_0_data_master_byteenable
	wire         mm_interconnect_0_cpu_0_jtag_debug_module_waitrequest;       // cpu_0:jtag_debug_module_waitrequest -> mm_interconnect_0:cpu_0_jtag_debug_module_waitrequest
	wire  [31:0] mm_interconnect_0_cpu_0_jtag_debug_module_writedata;         // mm_interconnect_0:cpu_0_jtag_debug_module_writedata -> cpu_0:jtag_debug_module_writedata
	wire   [8:0] mm_interconnect_0_cpu_0_jtag_debug_module_address;           // mm_interconnect_0:cpu_0_jtag_debug_module_address -> cpu_0:jtag_debug_module_address
	wire         mm_interconnect_0_cpu_0_jtag_debug_module_write;             // mm_interconnect_0:cpu_0_jtag_debug_module_write -> cpu_0:jtag_debug_module_write
	wire         mm_interconnect_0_cpu_0_jtag_debug_module_read;              // mm_interconnect_0:cpu_0_jtag_debug_module_read -> cpu_0:jtag_debug_module_read
	wire  [31:0] mm_interconnect_0_cpu_0_jtag_debug_module_readdata;          // cpu_0:jtag_debug_module_readdata -> mm_interconnect_0:cpu_0_jtag_debug_module_readdata
	wire         mm_interconnect_0_cpu_0_jtag_debug_module_debugaccess;       // mm_interconnect_0:cpu_0_jtag_debug_module_debugaccess -> cpu_0:jtag_debug_module_debugaccess
	wire   [3:0] mm_interconnect_0_cpu_0_jtag_debug_module_byteenable;        // mm_interconnect_0:cpu_0_jtag_debug_module_byteenable -> cpu_0:jtag_debug_module_byteenable
	wire         mm_interconnect_0_cpu_bridge_s0_waitrequest;                 // cpu_bridge:s0_waitrequest -> mm_interconnect_0:cpu_bridge_s0_waitrequest
	wire   [0:0] mm_interconnect_0_cpu_bridge_s0_burstcount;                  // mm_interconnect_0:cpu_bridge_s0_burstcount -> cpu_bridge:s0_burstcount
	wire  [31:0] mm_interconnect_0_cpu_bridge_s0_writedata;                   // mm_interconnect_0:cpu_bridge_s0_writedata -> cpu_bridge:s0_writedata
	wire  [21:0] mm_interconnect_0_cpu_bridge_s0_address;                     // mm_interconnect_0:cpu_bridge_s0_address -> cpu_bridge:s0_address
	wire         mm_interconnect_0_cpu_bridge_s0_write;                       // mm_interconnect_0:cpu_bridge_s0_write -> cpu_bridge:s0_write
	wire         mm_interconnect_0_cpu_bridge_s0_read;                        // mm_interconnect_0:cpu_bridge_s0_read -> cpu_bridge:s0_read
	wire  [31:0] mm_interconnect_0_cpu_bridge_s0_readdata;                    // cpu_bridge:s0_readdata -> mm_interconnect_0:cpu_bridge_s0_readdata
	wire         mm_interconnect_0_cpu_bridge_s0_debugaccess;                 // mm_interconnect_0:cpu_bridge_s0_debugaccess -> cpu_bridge:s0_debugaccess
	wire         mm_interconnect_0_cpu_bridge_s0_readdatavalid;               // cpu_bridge:s0_readdatavalid -> mm_interconnect_0:cpu_bridge_s0_readdatavalid
	wire   [3:0] mm_interconnect_0_cpu_bridge_s0_byteenable;                  // mm_interconnect_0:cpu_bridge_s0_byteenable -> cpu_bridge:s0_byteenable
	wire         mm_interconnect_0_flash_bridge_s0_waitrequest;               // flash_bridge:s0_waitrequest -> mm_interconnect_0:flash_bridge_s0_waitrequest
	wire   [0:0] mm_interconnect_0_flash_bridge_s0_burstcount;                // mm_interconnect_0:flash_bridge_s0_burstcount -> flash_bridge:s0_burstcount
	wire  [31:0] mm_interconnect_0_flash_bridge_s0_writedata;                 // mm_interconnect_0:flash_bridge_s0_writedata -> flash_bridge:s0_writedata
	wire  [21:0] mm_interconnect_0_flash_bridge_s0_address;                   // mm_interconnect_0:flash_bridge_s0_address -> flash_bridge:s0_address
	wire         mm_interconnect_0_flash_bridge_s0_write;                     // mm_interconnect_0:flash_bridge_s0_write -> flash_bridge:s0_write
	wire         mm_interconnect_0_flash_bridge_s0_read;                      // mm_interconnect_0:flash_bridge_s0_read -> flash_bridge:s0_read
	wire  [31:0] mm_interconnect_0_flash_bridge_s0_readdata;                  // flash_bridge:s0_readdata -> mm_interconnect_0:flash_bridge_s0_readdata
	wire         mm_interconnect_0_flash_bridge_s0_debugaccess;               // mm_interconnect_0:flash_bridge_s0_debugaccess -> flash_bridge:s0_debugaccess
	wire         mm_interconnect_0_flash_bridge_s0_readdatavalid;             // flash_bridge:s0_readdatavalid -> mm_interconnect_0:flash_bridge_s0_readdatavalid
	wire   [3:0] mm_interconnect_0_flash_bridge_s0_byteenable;                // mm_interconnect_0:flash_bridge_s0_byteenable -> flash_bridge:s0_byteenable
	wire         mm_interconnect_0_mm_bridge_0_s0_waitrequest;                // mm_bridge_0:s0_waitrequest -> mm_interconnect_0:mm_bridge_0_s0_waitrequest
	wire   [0:0] mm_interconnect_0_mm_bridge_0_s0_burstcount;                 // mm_interconnect_0:mm_bridge_0_s0_burstcount -> mm_bridge_0:s0_burstcount
	wire  [31:0] mm_interconnect_0_mm_bridge_0_s0_writedata;                  // mm_interconnect_0:mm_bridge_0_s0_writedata -> mm_bridge_0:s0_writedata
	wire  [19:0] mm_interconnect_0_mm_bridge_0_s0_address;                    // mm_interconnect_0:mm_bridge_0_s0_address -> mm_bridge_0:s0_address
	wire         mm_interconnect_0_mm_bridge_0_s0_write;                      // mm_interconnect_0:mm_bridge_0_s0_write -> mm_bridge_0:s0_write
	wire         mm_interconnect_0_mm_bridge_0_s0_read;                       // mm_interconnect_0:mm_bridge_0_s0_read -> mm_bridge_0:s0_read
	wire  [31:0] mm_interconnect_0_mm_bridge_0_s0_readdata;                   // mm_bridge_0:s0_readdata -> mm_interconnect_0:mm_bridge_0_s0_readdata
	wire         mm_interconnect_0_mm_bridge_0_s0_debugaccess;                // mm_interconnect_0:mm_bridge_0_s0_debugaccess -> mm_bridge_0:s0_debugaccess
	wire         mm_interconnect_0_mm_bridge_0_s0_readdatavalid;              // mm_bridge_0:s0_readdatavalid -> mm_interconnect_0:mm_bridge_0_s0_readdatavalid
	wire   [3:0] mm_interconnect_0_mm_bridge_0_s0_byteenable;                 // mm_interconnect_0:mm_bridge_0_s0_byteenable -> mm_bridge_0:s0_byteenable
	wire         cpu_0_tightly_coupled_instruction_master_0_waitrequest;      // mm_interconnect_1:cpu_0_tightly_coupled_instruction_master_0_waitrequest -> cpu_0:icm0_waitrequest
	wire  [27:0] cpu_0_tightly_coupled_instruction_master_0_address;          // cpu_0:icm0_address -> mm_interconnect_1:cpu_0_tightly_coupled_instruction_master_0_address
	wire         cpu_0_tightly_coupled_instruction_master_0_clken;            // cpu_0:icm0_clken -> mm_interconnect_1:cpu_0_tightly_coupled_instruction_master_0_clken
	wire         cpu_0_tightly_coupled_instruction_master_0_read;             // cpu_0:icm0_read -> mm_interconnect_1:cpu_0_tightly_coupled_instruction_master_0_read
	wire  [31:0] cpu_0_tightly_coupled_instruction_master_0_readdata;         // mm_interconnect_1:cpu_0_tightly_coupled_instruction_master_0_readdata -> cpu_0:icm0_readdata
	wire         cpu_0_tightly_coupled_instruction_master_0_readdatavalid;    // mm_interconnect_1:cpu_0_tightly_coupled_instruction_master_0_readdatavalid -> cpu_0:icm0_readdatavalid
	wire  [31:0] mm_interconnect_1_tc_mem_s1_writedata;                       // mm_interconnect_1:tc_mem_s1_writedata -> tc_mem:writedata
	wire  [12:0] mm_interconnect_1_tc_mem_s1_address;                         // mm_interconnect_1:tc_mem_s1_address -> tc_mem:address
	wire         mm_interconnect_1_tc_mem_s1_chipselect;                      // mm_interconnect_1:tc_mem_s1_chipselect -> tc_mem:chipselect
	wire         mm_interconnect_1_tc_mem_s1_clken;                           // mm_interconnect_1:tc_mem_s1_clken -> tc_mem:clken
	wire         mm_interconnect_1_tc_mem_s1_write;                           // mm_interconnect_1:tc_mem_s1_write -> tc_mem:write
	wire  [31:0] mm_interconnect_1_tc_mem_s1_readdata;                        // tc_mem:readdata -> mm_interconnect_1:tc_mem_s1_readdata
	wire   [3:0] mm_interconnect_1_tc_mem_s1_byteenable;                      // mm_interconnect_1:tc_mem_s1_byteenable -> tc_mem:byteenable
	wire         cpu_0_tightly_coupled_data_master_0_waitrequest;             // mm_interconnect_2:cpu_0_tightly_coupled_data_master_0_waitrequest -> cpu_0:dcm0_waitrequest
	wire  [31:0] cpu_0_tightly_coupled_data_master_0_writedata;               // cpu_0:dcm0_writedata -> mm_interconnect_2:cpu_0_tightly_coupled_data_master_0_writedata
	wire  [27:0] cpu_0_tightly_coupled_data_master_0_address;                 // cpu_0:dcm0_address -> mm_interconnect_2:cpu_0_tightly_coupled_data_master_0_address
	wire         cpu_0_tightly_coupled_data_master_0_clken;                   // cpu_0:dcm0_clken -> mm_interconnect_2:cpu_0_tightly_coupled_data_master_0_clken
	wire         cpu_0_tightly_coupled_data_master_0_write;                   // cpu_0:dcm0_write -> mm_interconnect_2:cpu_0_tightly_coupled_data_master_0_write
	wire         cpu_0_tightly_coupled_data_master_0_read;                    // cpu_0:dcm0_read -> mm_interconnect_2:cpu_0_tightly_coupled_data_master_0_read
	wire  [31:0] cpu_0_tightly_coupled_data_master_0_readdata;                // mm_interconnect_2:cpu_0_tightly_coupled_data_master_0_readdata -> cpu_0:dcm0_readdata
	wire   [3:0] cpu_0_tightly_coupled_data_master_0_byteenable;              // cpu_0:dcm0_byteenable -> mm_interconnect_2:cpu_0_tightly_coupled_data_master_0_byteenable
	wire         cpu_0_tightly_coupled_data_master_0_readdatavalid;           // mm_interconnect_2:cpu_0_tightly_coupled_data_master_0_readdatavalid -> cpu_0:dcm0_readdatavalid
	wire  [31:0] mm_interconnect_2_tc_mem_s2_writedata;                       // mm_interconnect_2:tc_mem_s2_writedata -> tc_mem:writedata2
	wire  [12:0] mm_interconnect_2_tc_mem_s2_address;                         // mm_interconnect_2:tc_mem_s2_address -> tc_mem:address2
	wire         mm_interconnect_2_tc_mem_s2_chipselect;                      // mm_interconnect_2:tc_mem_s2_chipselect -> tc_mem:chipselect2
	wire         mm_interconnect_2_tc_mem_s2_clken;                           // mm_interconnect_2:tc_mem_s2_clken -> tc_mem:clken2
	wire         mm_interconnect_2_tc_mem_s2_write;                           // mm_interconnect_2:tc_mem_s2_write -> tc_mem:write2
	wire  [31:0] mm_interconnect_2_tc_mem_s2_readdata;                        // tc_mem:readdata2 -> mm_interconnect_2:tc_mem_s2_readdata
	wire   [3:0] mm_interconnect_2_tc_mem_s2_byteenable;                      // mm_interconnect_2:tc_mem_s2_byteenable -> tc_mem:byteenable2
	wire   [0:0] mm_bridge_0_m0_burstcount;                                   // mm_bridge_0:m0_burstcount -> mm_interconnect_3:mm_bridge_0_m0_burstcount
	wire         mm_bridge_0_m0_waitrequest;                                  // mm_interconnect_3:mm_bridge_0_m0_waitrequest -> mm_bridge_0:m0_waitrequest
	wire  [19:0] mm_bridge_0_m0_address;                                      // mm_bridge_0:m0_address -> mm_interconnect_3:mm_bridge_0_m0_address
	wire  [31:0] mm_bridge_0_m0_writedata;                                    // mm_bridge_0:m0_writedata -> mm_interconnect_3:mm_bridge_0_m0_writedata
	wire         mm_bridge_0_m0_write;                                        // mm_bridge_0:m0_write -> mm_interconnect_3:mm_bridge_0_m0_write
	wire         mm_bridge_0_m0_read;                                         // mm_bridge_0:m0_read -> mm_interconnect_3:mm_bridge_0_m0_read
	wire  [31:0] mm_bridge_0_m0_readdata;                                     // mm_interconnect_3:mm_bridge_0_m0_readdata -> mm_bridge_0:m0_readdata
	wire         mm_bridge_0_m0_debugaccess;                                  // mm_bridge_0:m0_debugaccess -> mm_interconnect_3:mm_bridge_0_m0_debugaccess
	wire   [3:0] mm_bridge_0_m0_byteenable;                                   // mm_bridge_0:m0_byteenable -> mm_interconnect_3:mm_bridge_0_m0_byteenable
	wire         mm_bridge_0_m0_readdatavalid;                                // mm_interconnect_3:mm_bridge_0_m0_readdatavalid -> mm_bridge_0:m0_readdatavalid
	wire         mm_interconnect_3_jtag_uart_0_avalon_jtag_slave_waitrequest; // jtag_uart_0:av_waitrequest -> mm_interconnect_3:jtag_uart_0_avalon_jtag_slave_waitrequest
	wire  [31:0] mm_interconnect_3_jtag_uart_0_avalon_jtag_slave_writedata;   // mm_interconnect_3:jtag_uart_0_avalon_jtag_slave_writedata -> jtag_uart_0:av_writedata
	wire   [0:0] mm_interconnect_3_jtag_uart_0_avalon_jtag_slave_address;     // mm_interconnect_3:jtag_uart_0_avalon_jtag_slave_address -> jtag_uart_0:av_address
	wire         mm_interconnect_3_jtag_uart_0_avalon_jtag_slave_chipselect;  // mm_interconnect_3:jtag_uart_0_avalon_jtag_slave_chipselect -> jtag_uart_0:av_chipselect
	wire         mm_interconnect_3_jtag_uart_0_avalon_jtag_slave_write;       // mm_interconnect_3:jtag_uart_0_avalon_jtag_slave_write -> jtag_uart_0:av_write_n
	wire         mm_interconnect_3_jtag_uart_0_avalon_jtag_slave_read;        // mm_interconnect_3:jtag_uart_0_avalon_jtag_slave_read -> jtag_uart_0:av_read_n
	wire  [31:0] mm_interconnect_3_jtag_uart_0_avalon_jtag_slave_readdata;    // jtag_uart_0:av_readdata -> mm_interconnect_3:jtag_uart_0_avalon_jtag_slave_readdata
	wire         mm_interconnect_3_slow_bridge_s0_waitrequest;                // slow_bridge:s0_waitrequest -> mm_interconnect_3:slow_bridge_s0_waitrequest
	wire   [0:0] mm_interconnect_3_slow_bridge_s0_burstcount;                 // mm_interconnect_3:slow_bridge_s0_burstcount -> slow_bridge:s0_burstcount
	wire  [31:0] mm_interconnect_3_slow_bridge_s0_writedata;                  // mm_interconnect_3:slow_bridge_s0_writedata -> slow_bridge:s0_writedata
	wire  [18:0] mm_interconnect_3_slow_bridge_s0_address;                    // mm_interconnect_3:slow_bridge_s0_address -> slow_bridge:s0_address
	wire         mm_interconnect_3_slow_bridge_s0_write;                      // mm_interconnect_3:slow_bridge_s0_write -> slow_bridge:s0_write
	wire         mm_interconnect_3_slow_bridge_s0_read;                       // mm_interconnect_3:slow_bridge_s0_read -> slow_bridge:s0_read
	wire  [31:0] mm_interconnect_3_slow_bridge_s0_readdata;                   // slow_bridge:s0_readdata -> mm_interconnect_3:slow_bridge_s0_readdata
	wire         mm_interconnect_3_slow_bridge_s0_debugaccess;                // mm_interconnect_3:slow_bridge_s0_debugaccess -> slow_bridge:s0_debugaccess
	wire         mm_interconnect_3_slow_bridge_s0_readdatavalid;              // slow_bridge:s0_readdatavalid -> mm_interconnect_3:slow_bridge_s0_readdatavalid
	wire   [3:0] mm_interconnect_3_slow_bridge_s0_byteenable;                 // mm_interconnect_3:slow_bridge_s0_byteenable -> slow_bridge:s0_byteenable
	wire  [31:0] mm_interconnect_3_powerlink_led_s1_writedata;                // mm_interconnect_3:POWERLINK_LED_s1_writedata -> POWERLINK_LED:writedata
	wire   [2:0] mm_interconnect_3_powerlink_led_s1_address;                  // mm_interconnect_3:POWERLINK_LED_s1_address -> POWERLINK_LED:address
	wire         mm_interconnect_3_powerlink_led_s1_chipselect;               // mm_interconnect_3:POWERLINK_LED_s1_chipselect -> POWERLINK_LED:chipselect
	wire         mm_interconnect_3_powerlink_led_s1_write;                    // mm_interconnect_3:POWERLINK_LED_s1_write -> POWERLINK_LED:write_n
	wire  [31:0] mm_interconnect_3_powerlink_led_s1_readdata;                 // POWERLINK_LED:readdata -> mm_interconnect_3:POWERLINK_LED_s1_readdata
	wire  [31:0] mm_interconnect_3_benchmark_pio_s1_writedata;                // mm_interconnect_3:benchmark_pio_s1_writedata -> benchmark_pio:writedata
	wire   [2:0] mm_interconnect_3_benchmark_pio_s1_address;                  // mm_interconnect_3:benchmark_pio_s1_address -> benchmark_pio:address
	wire         mm_interconnect_3_benchmark_pio_s1_chipselect;               // mm_interconnect_3:benchmark_pio_s1_chipselect -> benchmark_pio:chipselect
	wire         mm_interconnect_3_benchmark_pio_s1_write;                    // mm_interconnect_3:benchmark_pio_s1_write -> benchmark_pio:write_n
	wire  [31:0] mm_interconnect_3_benchmark_pio_s1_readdata;                 // benchmark_pio:readdata -> mm_interconnect_3:benchmark_pio_s1_readdata
	wire  [15:0] mm_interconnect_3_timer_0_s1_writedata;                      // mm_interconnect_3:timer_0_s1_writedata -> timer_0:writedata
	wire   [2:0] mm_interconnect_3_timer_0_s1_address;                        // mm_interconnect_3:timer_0_s1_address -> timer_0:address
	wire         mm_interconnect_3_timer_0_s1_chipselect;                     // mm_interconnect_3:timer_0_s1_chipselect -> timer_0:chipselect
	wire         mm_interconnect_3_timer_0_s1_write;                          // mm_interconnect_3:timer_0_s1_write -> timer_0:write_n
	wire  [15:0] mm_interconnect_3_timer_0_s1_readdata;                       // timer_0:readdata -> mm_interconnect_3:timer_0_s1_readdata
	wire  [31:0] cpu_0_d_irq_irq;                                             // irq_mapper:sender_irq -> cpu_0:d_irq
	wire         irq_mapper_receiver0_irq;                                    // irq_synchronizer:sender_irq -> irq_mapper:receiver0_irq
	wire   [0:0] irq_synchronizer_receiver_irq;                               // timer_0:irq -> irq_synchronizer:receiver_irq
	wire         irq_mapper_receiver1_irq;                                    // irq_synchronizer_001:sender_irq -> irq_mapper:receiver1_irq
	wire   [0:0] irq_synchronizer_001_receiver_irq;                           // jtag_uart_0:av_irq -> irq_synchronizer_001:receiver_irq
	wire         irq_mapper_receiver2_irq;                                    // irq_synchronizer_002:sender_irq -> irq_mapper:receiver2_irq
	wire   [0:0] irq_synchronizer_002_receiver_irq;                           // sync_irq:sender0_irq -> irq_synchronizer_002:receiver_irq
	wire         irq_mapper_receiver3_irq;                                    // irq_synchronizer_003:sender_irq -> irq_mapper:receiver3_irq
	wire   [0:0] irq_synchronizer_003_receiver_irq;                           // mac_irq:sender0_irq -> irq_synchronizer_003:receiver_irq
	wire         irq_mapper_receiver4_irq;                                    // irq_synchronizer_004:sender_irq -> irq_mapper:receiver4_irq
	wire   [0:0] irq_synchronizer_004_receiver_irq;                           // gp_irq:sender0_irq -> irq_synchronizer_004:receiver_irq
	wire         irq_mapper_receiver5_irq;                                    // irq_synchronizer_005:sender_irq -> irq_mapper:receiver5_irq
	wire   [0:0] irq_synchronizer_005_receiver_irq;                           // gp_irq:sender1_irq -> irq_synchronizer_005:receiver_irq
	wire         irq_mapper_receiver6_irq;                                    // irq_synchronizer_006:sender_irq -> irq_mapper:receiver6_irq
	wire   [0:0] irq_synchronizer_006_receiver_irq;                           // gp_irq:sender2_irq -> irq_synchronizer_006:receiver_irq
	wire         irq_mapper_receiver7_irq;                                    // irq_synchronizer_007:sender_irq -> irq_mapper:receiver7_irq
	wire   [0:0] irq_synchronizer_007_receiver_irq;                           // gp_irq:sender3_irq -> irq_synchronizer_007:receiver_irq
	wire         rst_controller_reset_out_reset;                              // rst_controller:reset_out -> [cpu_0:reset_n, cpu_bridge:reset, irq_mapper:reset, irq_synchronizer:sender_reset, irq_synchronizer_001:sender_reset, irq_synchronizer_002:sender_reset, irq_synchronizer_003:sender_reset, irq_synchronizer_004:sender_reset, irq_synchronizer_005:sender_reset, irq_synchronizer_006:sender_reset, irq_synchronizer_007:sender_reset, mm_interconnect_0:cpu_0_reset_n_reset_bridge_in_reset_reset, mm_interconnect_1:cpu_0_reset_n_reset_bridge_in_reset_reset, mm_interconnect_2:cpu_0_reset_n_reset_bridge_in_reset_reset, rst_translator:in_reset, tc_mem:reset, tc_mem:reset2]
	wire         rst_controller_reset_out_reset_req;                          // rst_controller:reset_req -> [cpu_0:reset_req, rst_translator:reset_req_in, tc_mem:reset_req, tc_mem:reset_req2]
	wire         cpu_0_jtag_debug_module_reset_reset;                         // cpu_0:jtag_debug_module_resetrequest -> [rst_controller:reset_in1, rst_controller_001:reset_in2, rst_controller_002:reset_in0]
	wire         rst_controller_001_reset_out_reset;                          // rst_controller_001:reset_out -> [POWERLINK_LED:reset_n, benchmark_pio:reset_n, flash_bridge:reset, gp_irq:reset, irq_synchronizer:receiver_reset, irq_synchronizer_001:receiver_reset, jtag_uart_0:rst_n, mac_irq:reset, mm_bridge_0:reset, mm_interconnect_0:flash_bridge_reset_reset_bridge_in_reset_reset, mm_interconnect_3:mm_bridge_0_reset_reset_bridge_in_reset_reset, slow_bridge:reset, sync_irq:reset, timer_0:reset_n]

	soc_system_pcp_0_cpu_0 cpu_0 (
		.clk                                   (clk100_clk),                                               //                                  clk.clk
		.reset_n                               (~rst_controller_reset_out_reset),                          //                              reset_n.reset_n
		.reset_req                             (rst_controller_reset_out_reset_req),                       //                                     .reset_req
		.d_address                             (cpu_0_data_master_address),                                //                          data_master.address
		.d_byteenable                          (cpu_0_data_master_byteenable),                             //                                     .byteenable
		.d_read                                (cpu_0_data_master_read),                                   //                                     .read
		.d_readdata                            (cpu_0_data_master_readdata),                               //                                     .readdata
		.d_waitrequest                         (cpu_0_data_master_waitrequest),                            //                                     .waitrequest
		.d_write                               (cpu_0_data_master_write),                                  //                                     .write
		.d_writedata                           (cpu_0_data_master_writedata),                              //                                     .writedata
		.jtag_debug_module_debugaccess_to_roms (cpu_0_data_master_debugaccess),                            //                                     .debugaccess
		.i_address                             (cpu_0_instruction_master_address),                         //                   instruction_master.address
		.i_read                                (cpu_0_instruction_master_read),                            //                                     .read
		.i_readdata                            (cpu_0_instruction_master_readdata),                        //                                     .readdata
		.i_waitrequest                         (cpu_0_instruction_master_waitrequest),                     //                                     .waitrequest
		.i_readdatavalid                       (cpu_0_instruction_master_readdatavalid),                   //                                     .readdatavalid
		.dcm0_readdata                         (cpu_0_tightly_coupled_data_master_0_readdata),             //        tightly_coupled_data_master_0.readdata
		.dcm0_waitrequest                      (cpu_0_tightly_coupled_data_master_0_waitrequest),          //                                     .waitrequest
		.dcm0_readdatavalid                    (cpu_0_tightly_coupled_data_master_0_readdatavalid),        //                                     .readdatavalid
		.dcm0_address                          (cpu_0_tightly_coupled_data_master_0_address),              //                                     .address
		.dcm0_read                             (cpu_0_tightly_coupled_data_master_0_read),                 //                                     .read
		.dcm0_clken                            (cpu_0_tightly_coupled_data_master_0_clken),                //                                     .clken
		.dcm0_write                            (cpu_0_tightly_coupled_data_master_0_write),                //                                     .write
		.dcm0_writedata                        (cpu_0_tightly_coupled_data_master_0_writedata),            //                                     .writedata
		.dcm0_byteenable                       (cpu_0_tightly_coupled_data_master_0_byteenable),           //                                     .byteenable
		.icm0_readdata                         (cpu_0_tightly_coupled_instruction_master_0_readdata),      // tightly_coupled_instruction_master_0.readdata
		.icm0_waitrequest                      (cpu_0_tightly_coupled_instruction_master_0_waitrequest),   //                                     .waitrequest
		.icm0_readdatavalid                    (cpu_0_tightly_coupled_instruction_master_0_readdatavalid), //                                     .readdatavalid
		.icm0_address                          (cpu_0_tightly_coupled_instruction_master_0_address),       //                                     .address
		.icm0_read                             (cpu_0_tightly_coupled_instruction_master_0_read),          //                                     .read
		.icm0_clken                            (cpu_0_tightly_coupled_instruction_master_0_clken),         //                                     .clken
		.d_irq                                 (cpu_0_d_irq_irq),                                          //                                d_irq.irq
		.jtag_debug_module_resetrequest        (cpu_0_jtag_debug_module_reset_reset),                      //              jtag_debug_module_reset.reset
		.jtag_debug_module_address             (mm_interconnect_0_cpu_0_jtag_debug_module_address),        //                    jtag_debug_module.address
		.jtag_debug_module_byteenable          (mm_interconnect_0_cpu_0_jtag_debug_module_byteenable),     //                                     .byteenable
		.jtag_debug_module_debugaccess         (mm_interconnect_0_cpu_0_jtag_debug_module_debugaccess),    //                                     .debugaccess
		.jtag_debug_module_read                (mm_interconnect_0_cpu_0_jtag_debug_module_read),           //                                     .read
		.jtag_debug_module_readdata            (mm_interconnect_0_cpu_0_jtag_debug_module_readdata),       //                                     .readdata
		.jtag_debug_module_waitrequest         (mm_interconnect_0_cpu_0_jtag_debug_module_waitrequest),    //                                     .waitrequest
		.jtag_debug_module_write               (mm_interconnect_0_cpu_0_jtag_debug_module_write),          //                                     .write
		.jtag_debug_module_writedata           (mm_interconnect_0_cpu_0_jtag_debug_module_writedata),      //                                     .writedata
		.no_ci_readra                          (),                                                         //            custom_instruction_master.readra
		.cpu_resetrequest                      (cpu_resetrequest_resetrequest),                            //             cpu_resetrequest_conduit.export
		.cpu_resettaken                        (cpu_resetrequest_resettaken)                               //                                     .export
	);

	soc_system_pcp_0_tc_mem tc_mem (
		.clk         (clk100_clk),                             //   clk1.clk
		.address     (mm_interconnect_1_tc_mem_s1_address),    //     s1.address
		.clken       (mm_interconnect_1_tc_mem_s1_clken),      //       .clken
		.chipselect  (mm_interconnect_1_tc_mem_s1_chipselect), //       .chipselect
		.write       (mm_interconnect_1_tc_mem_s1_write),      //       .write
		.readdata    (mm_interconnect_1_tc_mem_s1_readdata),   //       .readdata
		.writedata   (mm_interconnect_1_tc_mem_s1_writedata),  //       .writedata
		.byteenable  (mm_interconnect_1_tc_mem_s1_byteenable), //       .byteenable
		.reset       (rst_controller_reset_out_reset),         // reset1.reset
		.reset_req   (rst_controller_reset_out_reset_req),     //       .reset_req
		.address2    (mm_interconnect_2_tc_mem_s2_address),    //     s2.address
		.chipselect2 (mm_interconnect_2_tc_mem_s2_chipselect), //       .chipselect
		.clken2      (mm_interconnect_2_tc_mem_s2_clken),      //       .clken
		.write2      (mm_interconnect_2_tc_mem_s2_write),      //       .write
		.readdata2   (mm_interconnect_2_tc_mem_s2_readdata),   //       .readdata
		.writedata2  (mm_interconnect_2_tc_mem_s2_writedata),  //       .writedata
		.byteenable2 (mm_interconnect_2_tc_mem_s2_byteenable), //       .byteenable
		.clk2        (clk100_clk),                             //   clk2.clk
		.reset2      (rst_controller_reset_out_reset),         // reset2.reset
		.reset_req2  (rst_controller_reset_out_reset_req)      //       .reset_req
	);

	soc_system_host_0_timer_0 timer_0 (
		.clk        (clk50_clk),                               //   clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),     // reset.reset_n
		.address    (mm_interconnect_3_timer_0_s1_address),    //    s1.address
		.writedata  (mm_interconnect_3_timer_0_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_3_timer_0_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_3_timer_0_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_3_timer_0_s1_write),     //      .write_n
		.irq        (irq_synchronizer_receiver_irq)            //   irq.irq
	);

	soc_system_pcp_0_benchmark_pio benchmark_pio (
		.clk        (clk50_clk),                                     //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),           //               reset.reset_n
		.address    (mm_interconnect_3_benchmark_pio_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_3_benchmark_pio_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_3_benchmark_pio_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_3_benchmark_pio_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_3_benchmark_pio_s1_readdata),   //                    .readdata
		.out_port   (benchmark_pio_external_connection_export)       // external_connection.export
	);

	soc_system_pcp_0_jtag_uart_0 jtag_uart_0 (
		.clk            (clk50_clk),                                                   //               clk.clk
		.rst_n          (~rst_controller_001_reset_out_reset),                         //             reset.reset_n
		.av_chipselect  (mm_interconnect_3_jtag_uart_0_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_3_jtag_uart_0_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_3_jtag_uart_0_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_3_jtag_uart_0_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_3_jtag_uart_0_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_3_jtag_uart_0_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_3_jtag_uart_0_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_synchronizer_001_receiver_irq)                            //               irq.irq
	);

	altera_avalon_mm_bridge #(
		.DATA_WIDTH        (32),
		.SYMBOL_WIDTH      (8),
		.HDL_ADDR_WIDTH    (19),
		.BURSTCOUNT_WIDTH  (1),
		.PIPELINE_COMMAND  (0),
		.PIPELINE_RESPONSE (0)
	) slow_bridge (
		.clk              (clk50_clk),                                      //   clk.clk
		.reset            (rst_controller_001_reset_out_reset),             // reset.reset
		.s0_waitrequest   (mm_interconnect_3_slow_bridge_s0_waitrequest),   //    s0.waitrequest
		.s0_readdata      (mm_interconnect_3_slow_bridge_s0_readdata),      //      .readdata
		.s0_readdatavalid (mm_interconnect_3_slow_bridge_s0_readdatavalid), //      .readdatavalid
		.s0_burstcount    (mm_interconnect_3_slow_bridge_s0_burstcount),    //      .burstcount
		.s0_writedata     (mm_interconnect_3_slow_bridge_s0_writedata),     //      .writedata
		.s0_address       (mm_interconnect_3_slow_bridge_s0_address),       //      .address
		.s0_write         (mm_interconnect_3_slow_bridge_s0_write),         //      .write
		.s0_read          (mm_interconnect_3_slow_bridge_s0_read),          //      .read
		.s0_byteenable    (mm_interconnect_3_slow_bridge_s0_byteenable),    //      .byteenable
		.s0_debugaccess   (mm_interconnect_3_slow_bridge_s0_debugaccess),   //      .debugaccess
		.m0_waitrequest   (slow_bridge_waitrequest),                        //    m0.waitrequest
		.m0_readdata      (slow_bridge_readdata),                           //      .readdata
		.m0_readdatavalid (slow_bridge_readdatavalid),                      //      .readdatavalid
		.m0_burstcount    (slow_bridge_burstcount),                         //      .burstcount
		.m0_writedata     (slow_bridge_writedata),                          //      .writedata
		.m0_address       (slow_bridge_address),                            //      .address
		.m0_write         (slow_bridge_write),                              //      .write
		.m0_read          (slow_bridge_read),                               //      .read
		.m0_byteenable    (slow_bridge_byteenable),                         //      .byteenable
		.m0_debugaccess   (slow_bridge_debugaccess)                         //      .debugaccess
	);

	altera_avalon_mm_bridge #(
		.DATA_WIDTH        (32),
		.SYMBOL_WIDTH      (8),
		.HDL_ADDR_WIDTH    (22),
		.BURSTCOUNT_WIDTH  (1),
		.PIPELINE_COMMAND  (0),
		.PIPELINE_RESPONSE (0)
	) cpu_bridge (
		.clk              (clk100_clk),                                    //   clk.clk
		.reset            (rst_controller_reset_out_reset),                // reset.reset
		.s0_waitrequest   (mm_interconnect_0_cpu_bridge_s0_waitrequest),   //    s0.waitrequest
		.s0_readdata      (mm_interconnect_0_cpu_bridge_s0_readdata),      //      .readdata
		.s0_readdatavalid (mm_interconnect_0_cpu_bridge_s0_readdatavalid), //      .readdatavalid
		.s0_burstcount    (mm_interconnect_0_cpu_bridge_s0_burstcount),    //      .burstcount
		.s0_writedata     (mm_interconnect_0_cpu_bridge_s0_writedata),     //      .writedata
		.s0_address       (mm_interconnect_0_cpu_bridge_s0_address),       //      .address
		.s0_write         (mm_interconnect_0_cpu_bridge_s0_write),         //      .write
		.s0_read          (mm_interconnect_0_cpu_bridge_s0_read),          //      .read
		.s0_byteenable    (mm_interconnect_0_cpu_bridge_s0_byteenable),    //      .byteenable
		.s0_debugaccess   (mm_interconnect_0_cpu_bridge_s0_debugaccess),   //      .debugaccess
		.m0_waitrequest   (cpu_bridge_waitrequest),                        //    m0.waitrequest
		.m0_readdata      (cpu_bridge_readdata),                           //      .readdata
		.m0_readdatavalid (cpu_bridge_readdatavalid),                      //      .readdatavalid
		.m0_burstcount    (cpu_bridge_burstcount),                         //      .burstcount
		.m0_writedata     (cpu_bridge_writedata),                          //      .writedata
		.m0_address       (cpu_bridge_address),                            //      .address
		.m0_write         (cpu_bridge_write),                              //      .write
		.m0_read          (cpu_bridge_read),                               //      .read
		.m0_byteenable    (cpu_bridge_byteenable),                         //      .byteenable
		.m0_debugaccess   (cpu_bridge_debugaccess)                         //      .debugaccess
	);

	altera_irq_bridge #(
		.IRQ_WIDTH (1)
	) sync_irq (
		.clk          (clk50_clk),                          //          clk.clk
		.receiver_irq (sync_irq_irq),                       // receiver_irq.irq
		.reset        (rst_controller_001_reset_out_reset), //    clk_reset.reset
		.sender0_irq  (irq_synchronizer_002_receiver_irq),  //  sender0_irq.irq
		.sender1_irq  (),                                   //  (terminated)
		.sender2_irq  (),                                   //  (terminated)
		.sender3_irq  (),                                   //  (terminated)
		.sender4_irq  (),                                   //  (terminated)
		.sender5_irq  (),                                   //  (terminated)
		.sender6_irq  (),                                   //  (terminated)
		.sender7_irq  (),                                   //  (terminated)
		.sender8_irq  (),                                   //  (terminated)
		.sender9_irq  (),                                   //  (terminated)
		.sender10_irq (),                                   //  (terminated)
		.sender11_irq (),                                   //  (terminated)
		.sender12_irq (),                                   //  (terminated)
		.sender13_irq (),                                   //  (terminated)
		.sender14_irq (),                                   //  (terminated)
		.sender15_irq (),                                   //  (terminated)
		.sender16_irq (),                                   //  (terminated)
		.sender17_irq (),                                   //  (terminated)
		.sender18_irq (),                                   //  (terminated)
		.sender19_irq (),                                   //  (terminated)
		.sender20_irq (),                                   //  (terminated)
		.sender21_irq (),                                   //  (terminated)
		.sender22_irq (),                                   //  (terminated)
		.sender23_irq (),                                   //  (terminated)
		.sender24_irq (),                                   //  (terminated)
		.sender25_irq (),                                   //  (terminated)
		.sender26_irq (),                                   //  (terminated)
		.sender27_irq (),                                   //  (terminated)
		.sender28_irq (),                                   //  (terminated)
		.sender29_irq (),                                   //  (terminated)
		.sender30_irq (),                                   //  (terminated)
		.sender31_irq ()                                    //  (terminated)
	);

	altera_irq_bridge #(
		.IRQ_WIDTH (1)
	) mac_irq (
		.clk          (clk50_clk),                          //          clk.clk
		.receiver_irq (mac_irq_irq),                        // receiver_irq.irq
		.reset        (rst_controller_001_reset_out_reset), //    clk_reset.reset
		.sender0_irq  (irq_synchronizer_003_receiver_irq),  //  sender0_irq.irq
		.sender1_irq  (),                                   //  (terminated)
		.sender2_irq  (),                                   //  (terminated)
		.sender3_irq  (),                                   //  (terminated)
		.sender4_irq  (),                                   //  (terminated)
		.sender5_irq  (),                                   //  (terminated)
		.sender6_irq  (),                                   //  (terminated)
		.sender7_irq  (),                                   //  (terminated)
		.sender8_irq  (),                                   //  (terminated)
		.sender9_irq  (),                                   //  (terminated)
		.sender10_irq (),                                   //  (terminated)
		.sender11_irq (),                                   //  (terminated)
		.sender12_irq (),                                   //  (terminated)
		.sender13_irq (),                                   //  (terminated)
		.sender14_irq (),                                   //  (terminated)
		.sender15_irq (),                                   //  (terminated)
		.sender16_irq (),                                   //  (terminated)
		.sender17_irq (),                                   //  (terminated)
		.sender18_irq (),                                   //  (terminated)
		.sender19_irq (),                                   //  (terminated)
		.sender20_irq (),                                   //  (terminated)
		.sender21_irq (),                                   //  (terminated)
		.sender22_irq (),                                   //  (terminated)
		.sender23_irq (),                                   //  (terminated)
		.sender24_irq (),                                   //  (terminated)
		.sender25_irq (),                                   //  (terminated)
		.sender26_irq (),                                   //  (terminated)
		.sender27_irq (),                                   //  (terminated)
		.sender28_irq (),                                   //  (terminated)
		.sender29_irq (),                                   //  (terminated)
		.sender30_irq (),                                   //  (terminated)
		.sender31_irq ()                                    //  (terminated)
	);

	altera_avalon_mm_bridge #(
		.DATA_WIDTH        (32),
		.SYMBOL_WIDTH      (8),
		.HDL_ADDR_WIDTH    (22),
		.BURSTCOUNT_WIDTH  (1),
		.PIPELINE_COMMAND  (0),
		.PIPELINE_RESPONSE (0)
	) flash_bridge (
		.clk              (clk50_clk),                                       //   clk.clk
		.reset            (rst_controller_001_reset_out_reset),              // reset.reset
		.s0_waitrequest   (mm_interconnect_0_flash_bridge_s0_waitrequest),   //    s0.waitrequest
		.s0_readdata      (mm_interconnect_0_flash_bridge_s0_readdata),      //      .readdata
		.s0_readdatavalid (mm_interconnect_0_flash_bridge_s0_readdatavalid), //      .readdatavalid
		.s0_burstcount    (mm_interconnect_0_flash_bridge_s0_burstcount),    //      .burstcount
		.s0_writedata     (mm_interconnect_0_flash_bridge_s0_writedata),     //      .writedata
		.s0_address       (mm_interconnect_0_flash_bridge_s0_address),       //      .address
		.s0_write         (mm_interconnect_0_flash_bridge_s0_write),         //      .write
		.s0_read          (mm_interconnect_0_flash_bridge_s0_read),          //      .read
		.s0_byteenable    (mm_interconnect_0_flash_bridge_s0_byteenable),    //      .byteenable
		.s0_debugaccess   (mm_interconnect_0_flash_bridge_s0_debugaccess),   //      .debugaccess
		.m0_waitrequest   (flash_bridge_waitrequest),                        //    m0.waitrequest
		.m0_readdata      (flash_bridge_readdata),                           //      .readdata
		.m0_readdatavalid (flash_bridge_readdatavalid),                      //      .readdatavalid
		.m0_burstcount    (flash_bridge_burstcount),                         //      .burstcount
		.m0_writedata     (flash_bridge_writedata),                          //      .writedata
		.m0_address       (flash_bridge_address),                            //      .address
		.m0_write         (flash_bridge_write),                              //      .write
		.m0_read          (flash_bridge_read),                               //      .read
		.m0_byteenable    (flash_bridge_byteenable),                         //      .byteenable
		.m0_debugaccess   (flash_bridge_debugaccess)                         //      .debugaccess
	);

	altera_irq_bridge #(
		.IRQ_WIDTH (4)
	) gp_irq (
		.clk          (clk50_clk),                          //          clk.clk
		.receiver_irq (gp_irq_irq),                         // receiver_irq.irq
		.reset        (rst_controller_001_reset_out_reset), //    clk_reset.reset
		.sender0_irq  (irq_synchronizer_004_receiver_irq),  //  sender0_irq.irq
		.sender1_irq  (irq_synchronizer_005_receiver_irq),  //  sender1_irq.irq
		.sender2_irq  (irq_synchronizer_006_receiver_irq),  //  sender2_irq.irq
		.sender3_irq  (irq_synchronizer_007_receiver_irq),  //  sender3_irq.irq
		.sender4_irq  (),                                   //  (terminated)
		.sender5_irq  (),                                   //  (terminated)
		.sender6_irq  (),                                   //  (terminated)
		.sender7_irq  (),                                   //  (terminated)
		.sender8_irq  (),                                   //  (terminated)
		.sender9_irq  (),                                   //  (terminated)
		.sender10_irq (),                                   //  (terminated)
		.sender11_irq (),                                   //  (terminated)
		.sender12_irq (),                                   //  (terminated)
		.sender13_irq (),                                   //  (terminated)
		.sender14_irq (),                                   //  (terminated)
		.sender15_irq (),                                   //  (terminated)
		.sender16_irq (),                                   //  (terminated)
		.sender17_irq (),                                   //  (terminated)
		.sender18_irq (),                                   //  (terminated)
		.sender19_irq (),                                   //  (terminated)
		.sender20_irq (),                                   //  (terminated)
		.sender21_irq (),                                   //  (terminated)
		.sender22_irq (),                                   //  (terminated)
		.sender23_irq (),                                   //  (terminated)
		.sender24_irq (),                                   //  (terminated)
		.sender25_irq (),                                   //  (terminated)
		.sender26_irq (),                                   //  (terminated)
		.sender27_irq (),                                   //  (terminated)
		.sender28_irq (),                                   //  (terminated)
		.sender29_irq (),                                   //  (terminated)
		.sender30_irq (),                                   //  (terminated)
		.sender31_irq ()                                    //  (terminated)
	);

	soc_system_pcp_0_POWERLINK_LED powerlink_led (
		.clk        (clk50_clk),                                     //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),           //               reset.reset_n
		.address    (mm_interconnect_3_powerlink_led_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_3_powerlink_led_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_3_powerlink_led_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_3_powerlink_led_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_3_powerlink_led_s1_readdata),   //                    .readdata
		.out_port   (powerlink_led_export)                           // external_connection.export
	);

	altera_avalon_mm_bridge #(
		.DATA_WIDTH        (32),
		.SYMBOL_WIDTH      (8),
		.HDL_ADDR_WIDTH    (20),
		.BURSTCOUNT_WIDTH  (1),
		.PIPELINE_COMMAND  (0),
		.PIPELINE_RESPONSE (0)
	) mm_bridge_0 (
		.clk              (clk50_clk),                                      //   clk.clk
		.reset            (rst_controller_001_reset_out_reset),             // reset.reset
		.s0_waitrequest   (mm_interconnect_0_mm_bridge_0_s0_waitrequest),   //    s0.waitrequest
		.s0_readdata      (mm_interconnect_0_mm_bridge_0_s0_readdata),      //      .readdata
		.s0_readdatavalid (mm_interconnect_0_mm_bridge_0_s0_readdatavalid), //      .readdatavalid
		.s0_burstcount    (mm_interconnect_0_mm_bridge_0_s0_burstcount),    //      .burstcount
		.s0_writedata     (mm_interconnect_0_mm_bridge_0_s0_writedata),     //      .writedata
		.s0_address       (mm_interconnect_0_mm_bridge_0_s0_address),       //      .address
		.s0_write         (mm_interconnect_0_mm_bridge_0_s0_write),         //      .write
		.s0_read          (mm_interconnect_0_mm_bridge_0_s0_read),          //      .read
		.s0_byteenable    (mm_interconnect_0_mm_bridge_0_s0_byteenable),    //      .byteenable
		.s0_debugaccess   (mm_interconnect_0_mm_bridge_0_s0_debugaccess),   //      .debugaccess
		.m0_waitrequest   (mm_bridge_0_m0_waitrequest),                     //    m0.waitrequest
		.m0_readdata      (mm_bridge_0_m0_readdata),                        //      .readdata
		.m0_readdatavalid (mm_bridge_0_m0_readdatavalid),                   //      .readdatavalid
		.m0_burstcount    (mm_bridge_0_m0_burstcount),                      //      .burstcount
		.m0_writedata     (mm_bridge_0_m0_writedata),                       //      .writedata
		.m0_address       (mm_bridge_0_m0_address),                         //      .address
		.m0_write         (mm_bridge_0_m0_write),                           //      .write
		.m0_read          (mm_bridge_0_m0_read),                            //      .read
		.m0_byteenable    (mm_bridge_0_m0_byteenable),                      //      .byteenable
		.m0_debugaccess   (mm_bridge_0_m0_debugaccess)                      //      .debugaccess
	);

	soc_system_pcp_0_mm_interconnect_0 mm_interconnect_0 (
		.clk100_clk_clk                                 (clk100_clk),                                            //                               clk100_clk.clk
		.clk50_clk_clk                                  (clk50_clk),                                             //                                clk50_clk.clk
		.cpu_0_reset_n_reset_bridge_in_reset_reset      (rst_controller_reset_out_reset),                        //      cpu_0_reset_n_reset_bridge_in_reset.reset
		.flash_bridge_reset_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),                    // flash_bridge_reset_reset_bridge_in_reset.reset
		.cpu_0_data_master_address                      (cpu_0_data_master_address),                             //                        cpu_0_data_master.address
		.cpu_0_data_master_waitrequest                  (cpu_0_data_master_waitrequest),                         //                                         .waitrequest
		.cpu_0_data_master_byteenable                   (cpu_0_data_master_byteenable),                          //                                         .byteenable
		.cpu_0_data_master_read                         (cpu_0_data_master_read),                                //                                         .read
		.cpu_0_data_master_readdata                     (cpu_0_data_master_readdata),                            //                                         .readdata
		.cpu_0_data_master_write                        (cpu_0_data_master_write),                               //                                         .write
		.cpu_0_data_master_writedata                    (cpu_0_data_master_writedata),                           //                                         .writedata
		.cpu_0_data_master_debugaccess                  (cpu_0_data_master_debugaccess),                         //                                         .debugaccess
		.cpu_0_instruction_master_address               (cpu_0_instruction_master_address),                      //                 cpu_0_instruction_master.address
		.cpu_0_instruction_master_waitrequest           (cpu_0_instruction_master_waitrequest),                  //                                         .waitrequest
		.cpu_0_instruction_master_read                  (cpu_0_instruction_master_read),                         //                                         .read
		.cpu_0_instruction_master_readdata              (cpu_0_instruction_master_readdata),                     //                                         .readdata
		.cpu_0_instruction_master_readdatavalid         (cpu_0_instruction_master_readdatavalid),                //                                         .readdatavalid
		.cpu_0_jtag_debug_module_address                (mm_interconnect_0_cpu_0_jtag_debug_module_address),     //                  cpu_0_jtag_debug_module.address
		.cpu_0_jtag_debug_module_write                  (mm_interconnect_0_cpu_0_jtag_debug_module_write),       //                                         .write
		.cpu_0_jtag_debug_module_read                   (mm_interconnect_0_cpu_0_jtag_debug_module_read),        //                                         .read
		.cpu_0_jtag_debug_module_readdata               (mm_interconnect_0_cpu_0_jtag_debug_module_readdata),    //                                         .readdata
		.cpu_0_jtag_debug_module_writedata              (mm_interconnect_0_cpu_0_jtag_debug_module_writedata),   //                                         .writedata
		.cpu_0_jtag_debug_module_byteenable             (mm_interconnect_0_cpu_0_jtag_debug_module_byteenable),  //                                         .byteenable
		.cpu_0_jtag_debug_module_waitrequest            (mm_interconnect_0_cpu_0_jtag_debug_module_waitrequest), //                                         .waitrequest
		.cpu_0_jtag_debug_module_debugaccess            (mm_interconnect_0_cpu_0_jtag_debug_module_debugaccess), //                                         .debugaccess
		.cpu_bridge_s0_address                          (mm_interconnect_0_cpu_bridge_s0_address),               //                            cpu_bridge_s0.address
		.cpu_bridge_s0_write                            (mm_interconnect_0_cpu_bridge_s0_write),                 //                                         .write
		.cpu_bridge_s0_read                             (mm_interconnect_0_cpu_bridge_s0_read),                  //                                         .read
		.cpu_bridge_s0_readdata                         (mm_interconnect_0_cpu_bridge_s0_readdata),              //                                         .readdata
		.cpu_bridge_s0_writedata                        (mm_interconnect_0_cpu_bridge_s0_writedata),             //                                         .writedata
		.cpu_bridge_s0_burstcount                       (mm_interconnect_0_cpu_bridge_s0_burstcount),            //                                         .burstcount
		.cpu_bridge_s0_byteenable                       (mm_interconnect_0_cpu_bridge_s0_byteenable),            //                                         .byteenable
		.cpu_bridge_s0_readdatavalid                    (mm_interconnect_0_cpu_bridge_s0_readdatavalid),         //                                         .readdatavalid
		.cpu_bridge_s0_waitrequest                      (mm_interconnect_0_cpu_bridge_s0_waitrequest),           //                                         .waitrequest
		.cpu_bridge_s0_debugaccess                      (mm_interconnect_0_cpu_bridge_s0_debugaccess),           //                                         .debugaccess
		.flash_bridge_s0_address                        (mm_interconnect_0_flash_bridge_s0_address),             //                          flash_bridge_s0.address
		.flash_bridge_s0_write                          (mm_interconnect_0_flash_bridge_s0_write),               //                                         .write
		.flash_bridge_s0_read                           (mm_interconnect_0_flash_bridge_s0_read),                //                                         .read
		.flash_bridge_s0_readdata                       (mm_interconnect_0_flash_bridge_s0_readdata),            //                                         .readdata
		.flash_bridge_s0_writedata                      (mm_interconnect_0_flash_bridge_s0_writedata),           //                                         .writedata
		.flash_bridge_s0_burstcount                     (mm_interconnect_0_flash_bridge_s0_burstcount),          //                                         .burstcount
		.flash_bridge_s0_byteenable                     (mm_interconnect_0_flash_bridge_s0_byteenable),          //                                         .byteenable
		.flash_bridge_s0_readdatavalid                  (mm_interconnect_0_flash_bridge_s0_readdatavalid),       //                                         .readdatavalid
		.flash_bridge_s0_waitrequest                    (mm_interconnect_0_flash_bridge_s0_waitrequest),         //                                         .waitrequest
		.flash_bridge_s0_debugaccess                    (mm_interconnect_0_flash_bridge_s0_debugaccess),         //                                         .debugaccess
		.mm_bridge_0_s0_address                         (mm_interconnect_0_mm_bridge_0_s0_address),              //                           mm_bridge_0_s0.address
		.mm_bridge_0_s0_write                           (mm_interconnect_0_mm_bridge_0_s0_write),                //                                         .write
		.mm_bridge_0_s0_read                            (mm_interconnect_0_mm_bridge_0_s0_read),                 //                                         .read
		.mm_bridge_0_s0_readdata                        (mm_interconnect_0_mm_bridge_0_s0_readdata),             //                                         .readdata
		.mm_bridge_0_s0_writedata                       (mm_interconnect_0_mm_bridge_0_s0_writedata),            //                                         .writedata
		.mm_bridge_0_s0_burstcount                      (mm_interconnect_0_mm_bridge_0_s0_burstcount),           //                                         .burstcount
		.mm_bridge_0_s0_byteenable                      (mm_interconnect_0_mm_bridge_0_s0_byteenable),           //                                         .byteenable
		.mm_bridge_0_s0_readdatavalid                   (mm_interconnect_0_mm_bridge_0_s0_readdatavalid),        //                                         .readdatavalid
		.mm_bridge_0_s0_waitrequest                     (mm_interconnect_0_mm_bridge_0_s0_waitrequest),          //                                         .waitrequest
		.mm_bridge_0_s0_debugaccess                     (mm_interconnect_0_mm_bridge_0_s0_debugaccess)           //                                         .debugaccess
	);

	soc_system_pcp_0_mm_interconnect_1 mm_interconnect_1 (
		.clk100_clk_clk                                           (clk100_clk),                                               //                                 clk100_clk.clk
		.cpu_0_reset_n_reset_bridge_in_reset_reset                (rst_controller_reset_out_reset),                           //        cpu_0_reset_n_reset_bridge_in_reset.reset
		.cpu_0_tightly_coupled_instruction_master_0_address       (cpu_0_tightly_coupled_instruction_master_0_address),       // cpu_0_tightly_coupled_instruction_master_0.address
		.cpu_0_tightly_coupled_instruction_master_0_waitrequest   (cpu_0_tightly_coupled_instruction_master_0_waitrequest),   //                                           .waitrequest
		.cpu_0_tightly_coupled_instruction_master_0_read          (cpu_0_tightly_coupled_instruction_master_0_read),          //                                           .read
		.cpu_0_tightly_coupled_instruction_master_0_readdata      (cpu_0_tightly_coupled_instruction_master_0_readdata),      //                                           .readdata
		.cpu_0_tightly_coupled_instruction_master_0_readdatavalid (cpu_0_tightly_coupled_instruction_master_0_readdatavalid), //                                           .readdatavalid
		.cpu_0_tightly_coupled_instruction_master_0_clken         (cpu_0_tightly_coupled_instruction_master_0_clken),         //                                           .clken
		.tc_mem_s1_address                                        (mm_interconnect_1_tc_mem_s1_address),                      //                                  tc_mem_s1.address
		.tc_mem_s1_write                                          (mm_interconnect_1_tc_mem_s1_write),                        //                                           .write
		.tc_mem_s1_readdata                                       (mm_interconnect_1_tc_mem_s1_readdata),                     //                                           .readdata
		.tc_mem_s1_writedata                                      (mm_interconnect_1_tc_mem_s1_writedata),                    //                                           .writedata
		.tc_mem_s1_byteenable                                     (mm_interconnect_1_tc_mem_s1_byteenable),                   //                                           .byteenable
		.tc_mem_s1_chipselect                                     (mm_interconnect_1_tc_mem_s1_chipselect),                   //                                           .chipselect
		.tc_mem_s1_clken                                          (mm_interconnect_1_tc_mem_s1_clken)                         //                                           .clken
	);

	soc_system_pcp_0_mm_interconnect_2 mm_interconnect_2 (
		.clk100_clk_clk                                    (clk100_clk),                                        //                          clk100_clk.clk
		.cpu_0_reset_n_reset_bridge_in_reset_reset         (rst_controller_reset_out_reset),                    // cpu_0_reset_n_reset_bridge_in_reset.reset
		.cpu_0_tightly_coupled_data_master_0_address       (cpu_0_tightly_coupled_data_master_0_address),       // cpu_0_tightly_coupled_data_master_0.address
		.cpu_0_tightly_coupled_data_master_0_waitrequest   (cpu_0_tightly_coupled_data_master_0_waitrequest),   //                                    .waitrequest
		.cpu_0_tightly_coupled_data_master_0_byteenable    (cpu_0_tightly_coupled_data_master_0_byteenable),    //                                    .byteenable
		.cpu_0_tightly_coupled_data_master_0_read          (cpu_0_tightly_coupled_data_master_0_read),          //                                    .read
		.cpu_0_tightly_coupled_data_master_0_readdata      (cpu_0_tightly_coupled_data_master_0_readdata),      //                                    .readdata
		.cpu_0_tightly_coupled_data_master_0_readdatavalid (cpu_0_tightly_coupled_data_master_0_readdatavalid), //                                    .readdatavalid
		.cpu_0_tightly_coupled_data_master_0_write         (cpu_0_tightly_coupled_data_master_0_write),         //                                    .write
		.cpu_0_tightly_coupled_data_master_0_writedata     (cpu_0_tightly_coupled_data_master_0_writedata),     //                                    .writedata
		.cpu_0_tightly_coupled_data_master_0_clken         (cpu_0_tightly_coupled_data_master_0_clken),         //                                    .clken
		.tc_mem_s2_address                                 (mm_interconnect_2_tc_mem_s2_address),               //                           tc_mem_s2.address
		.tc_mem_s2_write                                   (mm_interconnect_2_tc_mem_s2_write),                 //                                    .write
		.tc_mem_s2_readdata                                (mm_interconnect_2_tc_mem_s2_readdata),              //                                    .readdata
		.tc_mem_s2_writedata                               (mm_interconnect_2_tc_mem_s2_writedata),             //                                    .writedata
		.tc_mem_s2_byteenable                              (mm_interconnect_2_tc_mem_s2_byteenable),            //                                    .byteenable
		.tc_mem_s2_chipselect                              (mm_interconnect_2_tc_mem_s2_chipselect),            //                                    .chipselect
		.tc_mem_s2_clken                                   (mm_interconnect_2_tc_mem_s2_clken)                  //                                    .clken
	);

	soc_system_pcp_0_mm_interconnect_3 mm_interconnect_3 (
		.clk50_clk_clk                                 (clk50_clk),                                                   //                               clk50_clk.clk
		.mm_bridge_0_reset_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),                          // mm_bridge_0_reset_reset_bridge_in_reset.reset
		.mm_bridge_0_m0_address                        (mm_bridge_0_m0_address),                                      //                          mm_bridge_0_m0.address
		.mm_bridge_0_m0_waitrequest                    (mm_bridge_0_m0_waitrequest),                                  //                                        .waitrequest
		.mm_bridge_0_m0_burstcount                     (mm_bridge_0_m0_burstcount),                                   //                                        .burstcount
		.mm_bridge_0_m0_byteenable                     (mm_bridge_0_m0_byteenable),                                   //                                        .byteenable
		.mm_bridge_0_m0_read                           (mm_bridge_0_m0_read),                                         //                                        .read
		.mm_bridge_0_m0_readdata                       (mm_bridge_0_m0_readdata),                                     //                                        .readdata
		.mm_bridge_0_m0_readdatavalid                  (mm_bridge_0_m0_readdatavalid),                                //                                        .readdatavalid
		.mm_bridge_0_m0_write                          (mm_bridge_0_m0_write),                                        //                                        .write
		.mm_bridge_0_m0_writedata                      (mm_bridge_0_m0_writedata),                                    //                                        .writedata
		.mm_bridge_0_m0_debugaccess                    (mm_bridge_0_m0_debugaccess),                                  //                                        .debugaccess
		.benchmark_pio_s1_address                      (mm_interconnect_3_benchmark_pio_s1_address),                  //                        benchmark_pio_s1.address
		.benchmark_pio_s1_write                        (mm_interconnect_3_benchmark_pio_s1_write),                    //                                        .write
		.benchmark_pio_s1_readdata                     (mm_interconnect_3_benchmark_pio_s1_readdata),                 //                                        .readdata
		.benchmark_pio_s1_writedata                    (mm_interconnect_3_benchmark_pio_s1_writedata),                //                                        .writedata
		.benchmark_pio_s1_chipselect                   (mm_interconnect_3_benchmark_pio_s1_chipselect),               //                                        .chipselect
		.jtag_uart_0_avalon_jtag_slave_address         (mm_interconnect_3_jtag_uart_0_avalon_jtag_slave_address),     //           jtag_uart_0_avalon_jtag_slave.address
		.jtag_uart_0_avalon_jtag_slave_write           (mm_interconnect_3_jtag_uart_0_avalon_jtag_slave_write),       //                                        .write
		.jtag_uart_0_avalon_jtag_slave_read            (mm_interconnect_3_jtag_uart_0_avalon_jtag_slave_read),        //                                        .read
		.jtag_uart_0_avalon_jtag_slave_readdata        (mm_interconnect_3_jtag_uart_0_avalon_jtag_slave_readdata),    //                                        .readdata
		.jtag_uart_0_avalon_jtag_slave_writedata       (mm_interconnect_3_jtag_uart_0_avalon_jtag_slave_writedata),   //                                        .writedata
		.jtag_uart_0_avalon_jtag_slave_waitrequest     (mm_interconnect_3_jtag_uart_0_avalon_jtag_slave_waitrequest), //                                        .waitrequest
		.jtag_uart_0_avalon_jtag_slave_chipselect      (mm_interconnect_3_jtag_uart_0_avalon_jtag_slave_chipselect),  //                                        .chipselect
		.POWERLINK_LED_s1_address                      (mm_interconnect_3_powerlink_led_s1_address),                  //                        POWERLINK_LED_s1.address
		.POWERLINK_LED_s1_write                        (mm_interconnect_3_powerlink_led_s1_write),                    //                                        .write
		.POWERLINK_LED_s1_readdata                     (mm_interconnect_3_powerlink_led_s1_readdata),                 //                                        .readdata
		.POWERLINK_LED_s1_writedata                    (mm_interconnect_3_powerlink_led_s1_writedata),                //                                        .writedata
		.POWERLINK_LED_s1_chipselect                   (mm_interconnect_3_powerlink_led_s1_chipselect),               //                                        .chipselect
		.slow_bridge_s0_address                        (mm_interconnect_3_slow_bridge_s0_address),                    //                          slow_bridge_s0.address
		.slow_bridge_s0_write                          (mm_interconnect_3_slow_bridge_s0_write),                      //                                        .write
		.slow_bridge_s0_read                           (mm_interconnect_3_slow_bridge_s0_read),                       //                                        .read
		.slow_bridge_s0_readdata                       (mm_interconnect_3_slow_bridge_s0_readdata),                   //                                        .readdata
		.slow_bridge_s0_writedata                      (mm_interconnect_3_slow_bridge_s0_writedata),                  //                                        .writedata
		.slow_bridge_s0_burstcount                     (mm_interconnect_3_slow_bridge_s0_burstcount),                 //                                        .burstcount
		.slow_bridge_s0_byteenable                     (mm_interconnect_3_slow_bridge_s0_byteenable),                 //                                        .byteenable
		.slow_bridge_s0_readdatavalid                  (mm_interconnect_3_slow_bridge_s0_readdatavalid),              //                                        .readdatavalid
		.slow_bridge_s0_waitrequest                    (mm_interconnect_3_slow_bridge_s0_waitrequest),                //                                        .waitrequest
		.slow_bridge_s0_debugaccess                    (mm_interconnect_3_slow_bridge_s0_debugaccess),                //                                        .debugaccess
		.timer_0_s1_address                            (mm_interconnect_3_timer_0_s1_address),                        //                              timer_0_s1.address
		.timer_0_s1_write                              (mm_interconnect_3_timer_0_s1_write),                          //                                        .write
		.timer_0_s1_readdata                           (mm_interconnect_3_timer_0_s1_readdata),                       //                                        .readdata
		.timer_0_s1_writedata                          (mm_interconnect_3_timer_0_s1_writedata),                      //                                        .writedata
		.timer_0_s1_chipselect                         (mm_interconnect_3_timer_0_s1_chipselect)                      //                                        .chipselect
	);

	soc_system_pcp_0_irq_mapper irq_mapper (
		.clk           (clk100_clk),                     //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),       // receiver2.irq
		.receiver3_irq (irq_mapper_receiver3_irq),       // receiver3.irq
		.receiver4_irq (irq_mapper_receiver4_irq),       // receiver4.irq
		.receiver5_irq (irq_mapper_receiver5_irq),       // receiver5.irq
		.receiver6_irq (irq_mapper_receiver6_irq),       // receiver6.irq
		.receiver7_irq (irq_mapper_receiver7_irq),       // receiver7.irq
		.sender_irq    (cpu_0_d_irq_irq)                 //    sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer (
		.receiver_clk   (clk50_clk),                          //       receiver_clk.clk
		.sender_clk     (clk100_clk),                         //         sender_clk.clk
		.receiver_reset (rst_controller_001_reset_out_reset), // receiver_clk_reset.reset
		.sender_reset   (rst_controller_reset_out_reset),     //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_receiver_irq),      //           receiver.irq
		.sender_irq     (irq_mapper_receiver0_irq)            //             sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer_001 (
		.receiver_clk   (clk50_clk),                          //       receiver_clk.clk
		.sender_clk     (clk100_clk),                         //         sender_clk.clk
		.receiver_reset (rst_controller_001_reset_out_reset), // receiver_clk_reset.reset
		.sender_reset   (rst_controller_reset_out_reset),     //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_001_receiver_irq),  //           receiver.irq
		.sender_irq     (irq_mapper_receiver1_irq)            //             sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer_002 (
		.receiver_clk   (clk100_clk),                        //       receiver_clk.clk
		.sender_clk     (clk100_clk),                        //         sender_clk.clk
		.receiver_reset (),                                  // receiver_clk_reset.reset
		.sender_reset   (rst_controller_reset_out_reset),    //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_002_receiver_irq), //           receiver.irq
		.sender_irq     (irq_mapper_receiver2_irq)           //             sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer_003 (
		.receiver_clk   (clk100_clk),                        //       receiver_clk.clk
		.sender_clk     (clk100_clk),                        //         sender_clk.clk
		.receiver_reset (),                                  // receiver_clk_reset.reset
		.sender_reset   (rst_controller_reset_out_reset),    //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_003_receiver_irq), //           receiver.irq
		.sender_irq     (irq_mapper_receiver3_irq)           //             sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer_004 (
		.receiver_clk   (clk100_clk),                        //       receiver_clk.clk
		.sender_clk     (clk100_clk),                        //         sender_clk.clk
		.receiver_reset (),                                  // receiver_clk_reset.reset
		.sender_reset   (rst_controller_reset_out_reset),    //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_004_receiver_irq), //           receiver.irq
		.sender_irq     (irq_mapper_receiver4_irq)           //             sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer_005 (
		.receiver_clk   (clk100_clk),                        //       receiver_clk.clk
		.sender_clk     (clk100_clk),                        //         sender_clk.clk
		.receiver_reset (),                                  // receiver_clk_reset.reset
		.sender_reset   (rst_controller_reset_out_reset),    //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_005_receiver_irq), //           receiver.irq
		.sender_irq     (irq_mapper_receiver5_irq)           //             sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer_006 (
		.receiver_clk   (clk100_clk),                        //       receiver_clk.clk
		.sender_clk     (clk100_clk),                        //         sender_clk.clk
		.receiver_reset (),                                  // receiver_clk_reset.reset
		.sender_reset   (rst_controller_reset_out_reset),    //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_006_receiver_irq), //           receiver.irq
		.sender_irq     (irq_mapper_receiver6_irq)           //             sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer_007 (
		.receiver_clk   (clk100_clk),                        //       receiver_clk.clk
		.sender_clk     (clk100_clk),                        //         sender_clk.clk
		.receiver_reset (),                                  // receiver_clk_reset.reset
		.sender_reset   (rst_controller_reset_out_reset),    //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_007_receiver_irq), //           receiver.irq
		.sender_irq     (irq_mapper_receiver7_irq)           //             sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (3),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~rst_clk100_reset_n),                 // reset_in0.reset
		.reset_in1      (cpu_0_jtag_debug_module_reset_reset), // reset_in1.reset
		.reset_in2      (~rst_clk50_reset_n),                  // reset_in2.reset
		.clk            (clk100_clk),                          //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),      // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req),  //          .reset_req
		.reset_req_in0  (1'b0),                                // (terminated)
		.reset_req_in1  (1'b0),                                // (terminated)
		.reset_req_in2  (1'b0),                                // (terminated)
		.reset_in3      (1'b0),                                // (terminated)
		.reset_req_in3  (1'b0),                                // (terminated)
		.reset_in4      (1'b0),                                // (terminated)
		.reset_req_in4  (1'b0),                                // (terminated)
		.reset_in5      (1'b0),                                // (terminated)
		.reset_req_in5  (1'b0),                                // (terminated)
		.reset_in6      (1'b0),                                // (terminated)
		.reset_req_in6  (1'b0),                                // (terminated)
		.reset_in7      (1'b0),                                // (terminated)
		.reset_req_in7  (1'b0),                                // (terminated)
		.reset_in8      (1'b0),                                // (terminated)
		.reset_req_in8  (1'b0),                                // (terminated)
		.reset_in9      (1'b0),                                // (terminated)
		.reset_req_in9  (1'b0),                                // (terminated)
		.reset_in10     (1'b0),                                // (terminated)
		.reset_req_in10 (1'b0),                                // (terminated)
		.reset_in11     (1'b0),                                // (terminated)
		.reset_req_in11 (1'b0),                                // (terminated)
		.reset_in12     (1'b0),                                // (terminated)
		.reset_req_in12 (1'b0),                                // (terminated)
		.reset_in13     (1'b0),                                // (terminated)
		.reset_req_in13 (1'b0),                                // (terminated)
		.reset_in14     (1'b0),                                // (terminated)
		.reset_req_in14 (1'b0),                                // (terminated)
		.reset_in15     (1'b0),                                // (terminated)
		.reset_req_in15 (1'b0)                                 // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (3),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~rst_clk50_reset_n),                  // reset_in0.reset
		.reset_in1      (~rst_clk100_reset_n),                 // reset_in1.reset
		.reset_in2      (cpu_0_jtag_debug_module_reset_reset), // reset_in2.reset
		.clk            (clk50_clk),                           //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset),  // reset_out.reset
		.reset_req      (),                                    // (terminated)
		.reset_req_in0  (1'b0),                                // (terminated)
		.reset_req_in1  (1'b0),                                // (terminated)
		.reset_req_in2  (1'b0),                                // (terminated)
		.reset_in3      (1'b0),                                // (terminated)
		.reset_req_in3  (1'b0),                                // (terminated)
		.reset_in4      (1'b0),                                // (terminated)
		.reset_req_in4  (1'b0),                                // (terminated)
		.reset_in5      (1'b0),                                // (terminated)
		.reset_req_in5  (1'b0),                                // (terminated)
		.reset_in6      (1'b0),                                // (terminated)
		.reset_req_in6  (1'b0),                                // (terminated)
		.reset_in7      (1'b0),                                // (terminated)
		.reset_req_in7  (1'b0),                                // (terminated)
		.reset_in8      (1'b0),                                // (terminated)
		.reset_req_in8  (1'b0),                                // (terminated)
		.reset_in9      (1'b0),                                // (terminated)
		.reset_req_in9  (1'b0),                                // (terminated)
		.reset_in10     (1'b0),                                // (terminated)
		.reset_req_in10 (1'b0),                                // (terminated)
		.reset_in11     (1'b0),                                // (terminated)
		.reset_req_in11 (1'b0),                                // (terminated)
		.reset_in12     (1'b0),                                // (terminated)
		.reset_req_in12 (1'b0),                                // (terminated)
		.reset_in13     (1'b0),                                // (terminated)
		.reset_req_in13 (1'b0),                                // (terminated)
		.reset_in14     (1'b0),                                // (terminated)
		.reset_req_in14 (1'b0),                                // (terminated)
		.reset_in15     (1'b0),                                // (terminated)
		.reset_req_in15 (1'b0)                                 // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("both"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_002 (
		.reset_in0      (cpu_0_jtag_debug_module_reset_reset), // reset_in0.reset
		.clk            (clk100_clk),                          //       clk.clk
		.reset_out      (jtag_reset_reset),                    // reset_out.reset
		.reset_req      (),                                    // (terminated)
		.reset_req_in0  (1'b0),                                // (terminated)
		.reset_in1      (1'b0),                                // (terminated)
		.reset_req_in1  (1'b0),                                // (terminated)
		.reset_in2      (1'b0),                                // (terminated)
		.reset_req_in2  (1'b0),                                // (terminated)
		.reset_in3      (1'b0),                                // (terminated)
		.reset_req_in3  (1'b0),                                // (terminated)
		.reset_in4      (1'b0),                                // (terminated)
		.reset_req_in4  (1'b0),                                // (terminated)
		.reset_in5      (1'b0),                                // (terminated)
		.reset_req_in5  (1'b0),                                // (terminated)
		.reset_in6      (1'b0),                                // (terminated)
		.reset_req_in6  (1'b0),                                // (terminated)
		.reset_in7      (1'b0),                                // (terminated)
		.reset_req_in7  (1'b0),                                // (terminated)
		.reset_in8      (1'b0),                                // (terminated)
		.reset_req_in8  (1'b0),                                // (terminated)
		.reset_in9      (1'b0),                                // (terminated)
		.reset_req_in9  (1'b0),                                // (terminated)
		.reset_in10     (1'b0),                                // (terminated)
		.reset_req_in10 (1'b0),                                // (terminated)
		.reset_in11     (1'b0),                                // (terminated)
		.reset_req_in11 (1'b0),                                // (terminated)
		.reset_in12     (1'b0),                                // (terminated)
		.reset_req_in12 (1'b0),                                // (terminated)
		.reset_in13     (1'b0),                                // (terminated)
		.reset_req_in13 (1'b0),                                // (terminated)
		.reset_in14     (1'b0),                                // (terminated)
		.reset_req_in14 (1'b0),                                // (terminated)
		.reset_in15     (1'b0),                                // (terminated)
		.reset_req_in15 (1'b0)                                 // (terminated)
	);

endmodule
